module v (
	input [6:0] x,
	input [6:0] y,
	output reg [3:0] vga_r,
	output reg [3:0] vga_g,
	output reg [3:0] vga_b
);

	always @(*) begin
		if ((x == 7'd588 && y == 43) || (x == 482 && y == 7'd513) || (x == 7'd279 && y == 617) ||
		(x == 210 && y == 424) || (x == 7'd161 && y == 7'd596) || (x == 7'd356 && y == 503) ||
		(x == 290 && y == 7'd575) || (x == 7'd235 && y == 639) || (x == 7'd366 && y == 7'd42) ||
		(x == 7'd404 && y == 639) || (x == 599 && y == 238) || (x == 7'd632 && y == 7'd202) ||
		(x == 7'd185 && y == 7'd593) || (x == 7'd416 && y == 7'd448) || (x == 586 && y == 518) ||
		(x == 32 && y == 7'd272) || (x == 587 && y == 7'd415) || (x == 7'd394 && y == 419) ||
		(x == 518 && y == 213) || (x == 7'd17 && y == 7'd338) || (x == 7'd242 && y == 55) ||
		(x == 633 && y == 138) || (x == 7'd394 && y == 447) || (x == 487 && y == 7'd56) ||
		(x == 7'd554 && y == 7'd250) || (x == 199 && y == 630) || (x == 294 && y == 7'd572) ||
		(x == 281 && y == 7'd299) || (x == 534 && y == 324) || (x == 7'd459 && y == 7'd309) ||
		(x == 7'd275 && y == 7'd311) || (x == 12 && y == 7'd423) || (x == 68 && y == 7'd567) ||
		(x == 7'd4 && y == 332) || (x == 7'd199 && y == 481) || (x == 7'd17 && y == 7'd279) ||
		(x == 7'd482 && y == 80) || (x == 7'd7 && y == 151) || (x == 7'd599 && y == 7'd133) ||
		(x == 367 && y == 474) || (x == 522 && y == 459) || (x == 7'd323 && y == 296) ||
		(x == 7'd520 && y == 64) || (x == 7'd213 && y == 7'd49) || (x == 634 && y == 7'd200) ||
		(x == 143 && y == 7'd352) || (x == 489 && y == 509) || (x == 7'd380 && y == 7'd617) ||
		(x == 7'd415 && y == 120) || (x == 619 && y == 548) || (x == 7'd360 && y == 7'd461) ||
		(x == 367 && y == 486) || (x == 620 && y == 7'd15) || (x == 7'd458 && y == 362) ||
		(x == 7'd152 && y == 294) || (x == 412 && y == 514) || (x == 7'd165 && y == 160) ||
		(x == 7'd119 && y == 555) || (x == 306 && y == 445) || (x == 516 && y == 7'd635) ||
		(x == 562 && y == 145) || (x == 7'd459 && y == 239) || (x == 7'd508 && y == 7'd132) ||
		(x == 7'd305 && y == 7'd358) || (x == 546 && y == 7'd543) || (x == 7'd90 && y == 7'd137) ||
		(x == 7'd550 && y == 343) || (x == 488 && y == 583) || (x == 7'd558 && y == 476) ||
		(x == 504 && y == 7'd263) || (x == 7'd279 && y == 7'd516) || (x == 7'd631 && y == 7'd290) ||
		(x == 303 && y == 187) || (x == 328 && y == 150) || (x == 197 && y == 7'd635) ||
		(x == 379 && y == 7'd613) || (x == 449 && y == 445) || (x == 129 && y == 7'd570) ||
		(x == 7'd344 && y == 411) || (x == 520 && y == 7'd608) || (x == 7'd498 && y == 7'd424) ||
		(x == 458 && y == 7'd103) || (x == 454 && y == 7'd468) || (x == 7'd484 && y == 7'd399) ||
		(x == 265 && y == 7'd406) || (x == 7'd493 && y == 7'd541) || (x == 483 && y == 483) ||
		(x == 7'd486 && y == 7'd207) || (x == 269 && y == 483) || (x == 7'd154 && y == 7'd262) ||
		(x == 154 && y == 7'd256) || (x == 7'd613 && y == 7'd510) || (x == 7'd195 && y == 7'd394) ||
		(x == 346 && y == 7'd638) || (x == 7'd552 && y == 456) || (x == 7'd164 && y == 7'd412) ||
		(x == 7'd537 && y == 7'd310) || (x == 7'd370 && y == 7'd621) || (x == 7'd19 && y == 7'd84) ||
		(x == 7'd633 && y == 29) || (x == 7'd449 && y == 7'd617) || (x == 7'd119 && y == 7'd331) ||
		(x == 7'd147 && y == 7'd338) || (x == 474 && y == 7'd431) || (x == 349 && y == 275) ||
		(x == 7'd169 && y == 7'd489) || (x == 7'd617 && y == 7'd629) || (x == 7'd522 && y == 7'd364) ||
		(x == 556 && y == 255) || (x == 429 && y == 623) || (x == 7'd596 && y == 214) ||
		(x == 246 && y == 7'd215) || (x == 7'd566 && y == 7'd460) || (x == 538 && y == 424) ||
		(x == 465 && y == 7'd573) || (x == 7'd138 && y == 7'd556) || (x == 7'd318 && y == 7'd467) ||
		(x == 7'd82 && y == 7'd251) || (x == 409 && y == 233) || (x == 7'd573 && y == 56) ||
		(x == 7'd63 && y == 7'd219) || (x == 7'd190 && y == 7'd270) || (x == 7'd577 && y == 7'd81) ||
		(x == 426 && y == 7'd268) || (x == 380 && y == 7'd638) || (x == 435 && y == 7'd75) ||
		(x == 7'd211 && y == 213) || (x == 584 && y == 500) || (x == 493 && y == 229) ||
		(x == 174 && y == 529) || (x == 7'd418 && y == 7'd385) || (x == 637 && y == 7'd110) ||
		(x == 372 && y == 7'd50) || (x == 7'd439 && y == 7'd609) || (x == 109 && y == 7'd224) ||
		(x == 115 && y == 7'd547) || (x == 7'd99 && y == 318) || (x == 7'd579 && y == 51) ||
		(x == 7'd586 && y == 7'd254) || (x == 7'd594 && y == 169) || (x == 7'd111 && y == 7'd26) ||
		(x == 7'd353 && y == 511) || (x == 516 && y == 462) || (x == 547 && y == 7'd472) ||
		(x == 7'd211 && y == 7'd627) || (x == 7'd366 && y == 461) || (x == 386 && y == 284) ||
		(x == 7'd165 && y == 7'd368) || (x == 7'd431 && y == 459) || (x == 590 && y == 242) ||
		(x == 555 && y == 7'd637) || (x == 7'd608 && y == 7'd397) || (x == 199 && y == 7'd53) ||
		(x == 7'd412 && y == 565) || (x == 165 && y == 7'd388) || (x == 7'd486 && y == 7'd56) ||
		(x == 293 && y == 7'd120) || (x == 511 && y == 530) || (x == 7'd11 && y == 612) ||
		(x == 638 && y == 501) || (x == 263 && y == 509) || (x == 426 && y == 234) ||
		(x == 7'd374 && y == 7'd254) || (x == 7'd603 && y == 344) || (x == 7'd135 && y == 7'd606) ||
		(x == 7'd20 && y == 578) || (x == 7'd80 && y == 7'd339) || (x == 7'd581 && y == 7'd235) ||
		(x == 7'd249 && y == 180) || (x == 7'd92 && y == 228) || (x == 7'd620 && y == 407) ||
		(x == 7'd63 && y == 7'd244) || (x == 7'd230 && y == 7'd146) || (x == 7'd294 && y == 222) ||
		(x == 7'd323 && y == 474) || (x == 57 && y == 7'd454) || (x == 592 && y == 7'd96) ||
		(x == 7'd234 && y == 7'd225) || (x == 560 && y == 7'd635) || (x == 115 && y == 7'd309) ||
		(x == 7'd338 && y == 445) || (x == 311 && y == 7'd248) || (x == 251 && y == 7'd554) ||
		(x == 7'd22 && y == 518) || (x == 246 && y == 7'd2) || (x == 383 && y == 7'd386) ||
		(x == 7'd243 && y == 7'd397) || (x == 7'd275 && y == 7'd196) || (x == 545 && y == 7'd102) ||
		(x == 7'd47 && y == 589) || (x == 7'd5 && y == 7'd105) || (x == 7'd401 && y == 7'd276) ||
		(x == 7'd454 && y == 8) || (x == 69 && y == 7'd377) || (x == 392 && y == 420) ||
		(x == 7'd249 && y == 7'd411) || (x == 7'd98 && y == 350) || (x == 420 && y == 7'd609) ||
		(x == 7'd141 && y == 0) || (x == 195 && y == 7'd459) || (x == 443 && y == 505) ||
		(x == 209 && y == 7'd585) || (x == 7'd2 && y == 7'd453) || (x == 7'd605 && y == 7'd435) ||
		(x == 82 && y == 7'd580) || (x == 330 && y == 599) || (x == 315 && y == 412) ||
		(x == 7'd436 && y == 7'd567) || (x == 399 && y == 529) || (x == 7'd2 && y == 7'd50) ||
		(x == 344 && y == 7'd446) || (x == 7'd546 && y == 7'd191) || (x == 147 && y == 7'd417) ||
		(x == 326 && y == 7'd13) || (x == 7'd410 && y == 360) || (x == 7'd162 && y == 7'd371) ||
		(x == 401 && y == 219) || (x == 7'd135 && y == 7'd313) || (x == 188 && y == 274) ||
		(x == 387 && y == 7'd443) || (x == 256 && y == 7'd464) || (x == 402 && y == 7'd78) ||
		(x == 7'd411 && y == 273) || (x == 578 && y == 7'd356) || (x == 7'd185 && y == 7'd0) ||
		(x == 7'd233 && y == 7'd131) || (x == 7'd404 && y == 7'd308) || (x == 7'd389 && y == 12) ||
		(x == 429 && y == 618) || (x == 7'd556 && y == 219) || (x == 261 && y == 7'd478) ||
		(x == 7'd265 && y == 7'd222) || (x == 7'd341 && y == 7'd627) || (x == 421 && y == 7'd169) ||
		(x == 7'd622 && y == 7'd224) || (x == 7'd166 && y == 7'd245) || (x == 134 && y == 7'd317) ||
		(x == 340 && y == 259) || (x == 7'd234 && y == 7'd282) || (x == 7'd509 && y == 600) ||
		(x == 249 && y == 7'd522) || (x == 7'd406 && y == 7'd308) || (x == 7'd306 && y == 284) ||
		(x == 7'd444 && y == 7'd580) || (x == 7'd451 && y == 579) || (x == 7'd477 && y == 170) ||
		(x == 7'd317 && y == 7'd243) || (x == 148 && y == 625) || (x == 598 && y == 7'd118) ||
		(x == 101 && y == 7'd172) || (x == 212 && y == 606) || (x == 106 && y == 7'd226) ||
		(x == 489 && y == 7'd465) || (x == 255 && y == 7'd343) || (x == 7'd454 && y == 7'd584) ||
		(x == 7'd159 && y == 7'd67) || (x == 7'd447 && y == 7'd432) || (x == 7'd256 && y == 381) ||
		(x == 2 && y == 95) || (x == 7'd519 && y == 7'd194) || (x == 7'd403 && y == 7'd427) ||
		(x == 185 && y == 7'd15) || (x == 372 && y == 7'd394) || (x == 7'd82 && y == 7'd428) ||
		(x == 7'd216 && y == 346) || (x == 232 && y == 511) || (x == 7'd523 && y == 7'd246) ||
		(x == 625 && y == 7'd474) || (x == 137 && y == 483) || (x == 7'd185 && y == 440) ||
		(x == 7'd344 && y == 354) || (x == 7'd612 && y == 7'd166) || (x == 529 && y == 558) ||
		(x == 7'd192 && y == 7'd325) || (x == 7'd314 && y == 7'd619) || (x == 7'd636 && y == 7'd618) ||
		(x == 7'd12 && y == 572) || (x == 317 && y == 7'd177) || (x == 7'd603 && y == 238) ||
		(x == 7'd451 && y == 7'd245) || (x == 176 && y == 606) || (x == 190 && y == 7'd548) ||
		(x == 7'd242 && y == 586) || (x == 7'd478 && y == 7'd508) || (x == 7'd277 && y == 7'd412) ||
		(x == 477 && y == 294) || (x == 7'd636 && y == 570) || (x == 7'd46 && y == 7'd389) ||
		(x == 7'd603 && y == 606) || (x == 7'd152 && y == 7'd380) || (x == 7'd378 && y == 250) ||
		(x == 86 && y == 7'd425) || (x == 7'd465 && y == 7'd250) || (x == 7'd85 && y == 7'd215) ||
		(x == 7'd240 && y == 7'd159) || (x == 546 && y == 191) || (x == 406 && y == 7'd451) ||
		(x == 433 && y == 217) || (x == 7'd631 && y == 369) || (x == 7'd415 && y == 7'd210) ||
		(x == 456 && y == 346) || (x == 266 && y == 374) || (x == 377 && y == 211) ||
		(x == 404 && y == 498) || (x == 7'd301 && y == 184) || (x == 7'd455 && y == 7'd311) ||
		(x == 7'd585 && y == 233) || (x == 625 && y == 467) || (x == 140 && y == 7'd614) ||
		(x == 7'd290 && y == 7'd473) || (x == 7'd617 && y == 267) || (x == 7'd145 && y == 7'd550) ||
		(x == 220 && y == 509) || (x == 7'd323 && y == 191) || (x == 162 && y == 7'd72) ||
		(x == 7'd508 && y == 217) || (x == 589 && y == 7'd167) || (x == 584 && y == 7'd455) ||
		(x == 435 && y == 418) || (x == 7'd190 && y == 7'd143) || (x == 7'd419 && y == 160) ||
		(x == 572 && y == 567) || (x == 7'd450 && y == 7'd7) || (x == 539 && y == 7'd546) ||
		(x == 7'd225 && y == 7'd273) || (x == 7'd53 && y == 410) || (x == 7'd324 && y == 7'd519) ||
		(x == 7'd412 && y == 7'd36) || (x == 44 && y == 7'd233) || (x == 196 && y == 526) ||
		(x == 627 && y == 7'd429) || (x == 165 && y == 7'd445) || (x == 161 && y == 7'd532) ||
		(x == 7'd198 && y == 7'd626) || (x == 7'd479 && y == 7'd636) || (x == 7'd538 && y == 7'd157) ||
		(x == 7'd613 && y == 7'd634) || (x == 7'd110 && y == 466) || (x == 480 && y == 588) ||
		(x == 7'd265 && y == 7'd220) || (x == 7'd471 && y == 7'd242) || (x == 7'd282 && y == 334) ||
		(x == 7'd215 && y == 578) || (x == 7'd627 && y == 7'd190) || (x == 7'd374 && y == 634) ||
		(x == 495 && y == 7'd296) || (x == 7'd550 && y == 235) || (x == 112 && y == 112) ||
		(x == 251 && y == 461) || (x == 158 && y == 269) || (x == 397 && y == 7'd209) ||
		(x == 7'd194 && y == 7'd377) || (x == 178 && y == 430) || (x == 359 && y == 504) ||
		(x == 7'd335 && y == 7'd363) || (x == 7'd201 && y == 577) || (x == 399 && y == 473) ||
		(x == 561 && y == 190) || (x == 384 && y == 7'd488) || (x == 7'd275 && y == 7'd284) ||
		(x == 227 && y == 7'd612) || (x == 289 && y == 7'd326) || (x == 7'd477 && y == 227) ||
		(x == 7'd467 && y == 7'd473) || (x == 7'd94 && y == 515) || (x == 383 && y == 7'd572) ||
		(x == 467 && y == 306) || (x == 635 && y == 147) || (x == 592 && y == 407) ||
		(x == 590 && y == 213) || (x == 447 && y == 7'd64) || (x == 8 && y == 7'd332) ||
		(x == 400 && y == 7'd573) || (x == 222 && y == 220) || (x == 7'd371 && y == 7'd602) ||
		(x == 7'd108 && y == 96) || (x == 7'd572 && y == 7'd173) || (x == 451 && y == 543) ||
		(x == 7'd466 && y == 7'd385) || (x == 258 && y == 7'd299) || (x == 267 && y == 7'd186) ||
		(x == 7'd350 && y == 546) || (x == 7'd531 && y == 7'd464) || (x == 7'd143 && y == 7'd195) ||
		(x == 237 && y == 617) || (x == 399 && y == 542) || (x == 406 && y == 227) ||
		(x == 7'd224 && y == 11) || (x == 33 && y == 7'd617) || (x == 462 && y == 7'd402) ||
		(x == 373 && y == 226) || (x == 431 && y == 7'd512) || (x == 7'd149 && y == 7'd397) ||
		(x == 7'd374 && y == 7'd484) || (x == 7'd177 && y == 7'd446) || (x == 486 && y == 340) ||
		(x == 7'd373 && y == 7'd332) || (x == 570 && y == 502) || (x == 157 && y == 627) ||
		(x == 484 && y == 333) || (x == 24 && y == 7'd381) || (x == 7'd54 && y == 344) ||
		(x == 346 && y == 7'd397) || (x == 7'd525 && y == 7'd21) || (x == 7'd288 && y == 7'd165) ||
		(x == 7'd157 && y == 121) || (x == 7'd490 && y == 7'd506) || (x == 7'd564 && y == 7'd18) ||
		(x == 7'd36 && y == 289) || (x == 7'd181 && y == 547) || (x == 7'd498 && y == 7'd625) ||
		(x == 88 && y == 7'd379) || (x == 153 && y == 449) || (x == 7'd640 && y == 202) ||
		(x == 7'd157 && y == 7'd635) || (x == 558 && y == 550) || (x == 485 && y == 640) ||
		(x == 7'd540 && y == 7'd379) || (x == 348 && y == 7'd128) || (x == 26 && y == 7'd71) ||
		(x == 173 && y == 7'd557) || (x == 548 && y == 390) || (x == 7'd18 && y == 606) ||
		(x == 7'd382 && y == 429) || (x == 536 && y == 161) || (x == 485 && y == 262) ||
		(x == 7'd194 && y == 7'd318) || (x == 7'd494 && y == 7'd216) || (x == 7'd193 && y == 195) ||
		(x == 560 && y == 213) || (x == 7'd477 && y == 7'd637) || (x == 7'd167 && y == 185) ||
		(x == 267 && y == 7'd334) || (x == 7'd247 && y == 7'd394) || (x == 7'd24 && y == 324) ||
		(x == 7'd480 && y == 392) || (x == 2 && y == 124) || (x == 7'd550 && y == 27) ||
		(x == 7'd369 && y == 203) || (x == 7'd440 && y == 7'd341) || (x == 242 && y == 231) ||
		(x == 7'd517 && y == 267) || (x == 270 && y == 392) || (x == 316 && y == 7'd248) ||
		(x == 298 && y == 557) || (x == 181 && y == 443) || (x == 529 && y == 584) ||
		(x == 7'd506 && y == 7'd488) || (x == 7'd628 && y == 494) || (x == 240 && y == 294) ||
		(x == 7'd194 && y == 573) || (x == 7'd503 && y == 7'd163) || (x == 636 && y == 7'd165) ||
		(x == 7'd194 && y == 145) || (x == 7'd172 && y == 521) || (x == 59 && y == 7'd377) ||
		(x == 451 && y == 7'd355) || (x == 7'd327 && y == 7'd551) || (x == 7'd397 && y == 7'd341) ||
		(x == 7'd336 && y == 7'd509) || (x == 7'd189 && y == 7'd168) || (x == 7'd515 && y == 124) ||
		(x == 7'd127 && y == 357) || (x == 7'd165 && y == 7'd218) || (x == 7'd226 && y == 606) ||
		(x == 350 && y == 7'd435) || (x == 182 && y == 280) || (x == 424 && y == 219) ||
		(x == 7'd90 && y == 14) || (x == 7'd589 && y == 7'd155) || (x == 7'd494 && y == 7'd453) ||
		(x == 7'd320 && y == 61) || (x == 162 && y == 558) || (x == 220 && y == 630) ||
		(x == 176 && y == 574) || (x == 93 && y == 7'd270) || (x == 485 && y == 7'd405) ||
		(x == 7'd15 && y == 7'd292) || (x == 7'd154 && y == 249) || (x == 363 && y == 312) ||
		(x == 298 && y == 293) || (x == 465 && y == 7'd535) || (x == 475 && y == 7'd194) ||
		(x == 7'd120 && y == 346) || (x == 7'd155 && y == 7'd14) || (x == 7'd555 && y == 37) ||
		(x == 491 && y == 7'd609) || (x == 7'd237 && y == 7'd347) || (x == 7'd72 && y == 7'd1) ||
		(x == 7'd301 && y == 404) || (x == 7'd556 && y == 160) || (x == 511 && y == 300) ||
		(x == 7'd383 && y == 7'd530) || (x == 179 && y == 7'd464) || (x == 7'd244 && y == 151) ||
		(x == 7'd345 && y == 403) || (x == 536 && y == 7'd478) || (x == 554 && y == 629) ||
		(x == 247 && y == 216) || (x == 437 && y == 7'd596) || (x == 523 && y == 7'd388) ||
		(x == 7'd632 && y == 7'd466) || (x == 7'd271 && y == 7'd449) || (x == 343 && y == 7'd167) ||
		(x == 523 && y == 585) || (x == 425 && y == 307) || (x == 590 && y == 587) ||
		(x == 416 && y == 7'd250) || (x == 324 && y == 7'd66) || (x == 207 && y == 306) ||
		(x == 7'd567 && y == 7'd317) || (x == 7'd536 && y == 7'd309) || (x == 7'd174 && y == 568) ||
		(x == 127 && y == 7'd246) || (x == 445 && y == 7'd100) || (x == 170 && y == 7'd496) ||
		(x == 7'd194 && y == 7'd361) || (x == 617 && y == 7'd360) || (x == 7'd48 && y == 7'd14) ||
		(x == 7'd200 && y == 7'd78) || (x == 7'd341 && y == 325) || (x == 196 && y == 7'd12) ||
		(x == 7'd608 && y == 7'd566) || (x == 7'd136 && y == 532) || (x == 610 && y == 222) ||
		(x == 7'd32 && y == 7'd285) || (x == 7'd134 && y == 7'd263) || (x == 7'd499 && y == 7'd319) ||
		(x == 275 && y == 557) || (x == 7'd217 && y == 7'd614) || (x == 7'd515 && y == 7'd157) ||
		(x == 7'd356 && y == 7'd156) || (x == 199 && y == 7'd359) || (x == 515 && y == 224) ||
		(x == 7'd532 && y == 7'd503) || (x == 7'd426 && y == 7'd574) || (x == 496 && y == 7'd457) ||
		(x == 7'd631 && y == 7'd541) || (x == 7'd638 && y == 7'd556) || (x == 7'd230 && y == 488) ||
		(x == 7'd184 && y == 7'd210) || (x == 7'd448 && y == 7'd40) || (x == 580 && y == 156) ||
		(x == 268 && y == 470) || (x == 300 && y == 636) || (x == 7'd441 && y == 7'd637) ||
		(x == 7'd122 && y == 491) || (x == 125 && y == 52) || (x == 7'd617 && y == 7'd560) ||
		(x == 7'd499 && y == 162) || (x == 7'd113 && y == 512) || (x == 7'd486 && y == 7'd563) ||
		(x == 7'd71 && y == 7'd37) || (x == 323 && y == 157) || (x == 287 && y == 7'd32) ||
		(x == 7'd367 && y == 187) || (x == 7'd375 && y == 478) || (x == 495 && y == 620) ||
		(x == 7'd195 && y == 7'd180) || (x == 240 && y == 7'd41) || (x == 351 && y == 254) ||
		(x == 7'd584 && y == 7'd3) || (x == 7'd580 && y == 560) || (x == 7'd188 && y == 41) ||
		(x == 7'd517 && y == 7'd458) || (x == 7'd416 && y == 185) || (x == 124 && y == 7'd595) ||
		(x == 277 && y == 7'd423) || (x == 7'd158 && y == 7'd204) || (x == 7'd444 && y == 118) ||
		(x == 365 && y == 7'd104) || (x == 7'd412 && y == 7'd209) || (x == 7'd230 && y == 7'd229) ||
		(x == 7'd362 && y == 7'd539) || (x == 506 && y == 7'd515) || (x == 635 && y == 7'd67) ||
		(x == 7'd442 && y == 312) || (x == 7'd175 && y == 107) || (x == 7'd607 && y == 405) ||
		(x == 7'd532 && y == 7'd513) || (x == 7'd273 && y == 7'd139) || (x == 362 && y == 7'd15) ||
		(x == 7'd630 && y == 7'd419) || (x == 7'd21 && y == 7'd301) || (x == 7'd427 && y == 7'd239) ||
		(x == 256 && y == 7'd139) || (x == 7'd581 && y == 7'd494) || (x == 7'd131 && y == 7'd233) ||
		(x == 176 && y == 7'd307) || (x == 7'd426 && y == 7'd210) || (x == 291 && y == 7'd88) ||
		(x == 7'd236 && y == 7'd180) || (x == 456 && y == 7'd460) || (x == 622 && y == 228) ||
		(x == 529 && y == 496) || (x == 7'd333 && y == 7'd210) || (x == 437 && y == 7'd375) ||
		(x == 154 && y == 529) || (x == 7'd31 && y == 610) || (x == 165 && y == 459) ||
		(x == 7'd68 && y == 7'd210) || (x == 7'd59 && y == 149) || (x == 7'd119 && y == 386) ||
		(x == 7'd478 && y == 393) || (x == 7'd505 && y == 7'd122) || (x == 7'd254 && y == 7'd619) ||
		(x == 7'd377 && y == 153) || (x == 365 && y == 489) || (x == 268 && y == 305) ||
		(x == 7'd485 && y == 7'd467) || (x == 7'd358 && y == 7'd483) || (x == 282 && y == 140) ||
		(x == 7'd195 && y == 5) || (x == 168 && y == 285) || (x == 7'd550 && y == 7'd624) ||
		(x == 439 && y == 344) || (x == 433 && y == 7'd620) || (x == 7'd192 && y == 7'd115) ||
		(x == 7'd614 && y == 7'd487) || (x == 7'd29 && y == 7'd506) || (x == 610 && y == 7'd593) ||
		(x == 7'd293 && y == 7'd481) || (x == 7'd624 && y == 130) || (x == 7'd394 && y == 7'd472) ||
		(x == 221 && y == 312) || (x == 7'd328 && y == 594) || (x == 7'd371 && y == 7'd621) ||
		(x == 7'd622 && y == 550) || (x == 7'd397 && y == 7'd447) || (x == 7'd98 && y == 234) ||
		(x == 113 && y == 114) || (x == 337 && y == 7'd582) || (x == 7'd216 && y == 7'd270) ||
		(x == 217 && y == 517) || (x == 7'd359 && y == 7'd334) || (x == 566 && y == 7'd9) ||
		(x == 7'd336 && y == 102) || (x == 219 && y == 175) || (x == 7'd319 && y == 7'd447) ||
		(x == 7'd70 && y == 7'd123) || (x == 7'd147 && y == 7'd181) || (x == 172 && y == 221) ||
		(x == 7'd538 && y == 7'd520) || (x == 7'd197 && y == 143) || (x == 7'd488 && y == 7'd557) ||
		(x == 7'd159 && y == 7'd283) || (x == 7'd313 && y == 7'd325) || (x == 197 && y == 202) ||
		(x == 7'd622 && y == 349) || (x == 7'd495 && y == 7'd250) || (x == 412 && y == 326) ||
		(x == 7'd259 && y == 588) || (x == 7'd167 && y == 7'd107) || (x == 7'd475 && y == 7'd638) ||
		(x == 7'd383 && y == 7'd224) || (x == 538 && y == 350) || (x == 332 && y == 415) ||
		(x == 391 && y == 7'd128) || (x == 7'd254 && y == 310) || (x == 7'd534 && y == 532) ||
		(x == 7'd100 && y == 7'd205) || (x == 7'd304 && y == 164) || (x == 373 && y == 7'd451) ||
		(x == 483 && y == 7'd336) || (x == 7'd249 && y == 7'd260) || (x == 7'd515 && y == 7'd283) ||
		(x == 277 && y == 7'd265) || (x == 7'd319 && y == 7'd138) || (x == 290 && y == 7'd395) ||
		(x == 331 && y == 312) || (x == 622 && y == 306) || (x == 7'd138 && y == 370) ||
		(x == 146 && y == 631) || (x == 293 && y == 425) || (x == 582 && y == 573) ||
		(x == 504 && y == 7'd439) || (x == 7'd311 && y == 7'd552) || (x == 7'd19 && y == 7'd548) ||
		(x == 570 && y == 7'd307) || (x == 394 && y == 7'd49) || (x == 7'd361 && y == 130) ||
		(x == 366 && y == 7'd360) || (x == 473 && y == 7'd125) || (x == 7'd196 && y == 531) ||
		(x == 7'd567 && y == 7'd366) || (x == 7'd555 && y == 7'd9) || (x == 207 && y == 316) ||
		(x == 7'd628 && y == 7'd137) || (x == 7'd518 && y == 7'd526) || (x == 167 && y == 527) ||
		(x == 135 && y == 7'd21) || (x == 7'd372 && y == 7'd319) || (x == 7'd612 && y == 7'd230) ||
		(x == 7'd532 && y == 7'd583) || (x == 626 && y == 270) || (x == 7'd440 && y == 7'd531) ||
		(x == 7'd614 && y == 7'd298) || (x == 308 && y == 7'd278) || (x == 7'd599 && y == 130) ||
		(x == 7'd621 && y == 142) || (x == 7'd270 && y == 7'd190) || (x == 378 && y == 7'd26) ||
		(x == 7'd527 && y == 7'd297) || (x == 7'd31 && y == 262) || (x == 7'd392 && y == 446) ||
		(x == 500 && y == 200) || (x == 234 && y == 7'd296) || (x == 187 && y == 611) ||
		(x == 7'd244 && y == 7'd139) || (x == 7'd139 && y == 267) || (x == 543 && y == 454) ||
		(x == 7'd203 && y == 7'd385) || (x == 170 && y == 225) || (x == 7'd292 && y == 0) ||
		(x == 7'd215 && y == 465) || (x == 199 && y == 7'd90) || (x == 7'd619 && y == 7'd562) ||
		(x == 7'd412 && y == 7'd47) || (x == 361 && y == 326) || (x == 520 && y == 625) ||
		(x == 7'd376 && y == 7'd126) || (x == 7'd283 && y == 556) || (x == 622 && y == 191) ||
		(x == 7'd202 && y == 234) || (x == 7'd174 && y == 7'd619) || (x == 7'd346 && y == 7'd294) ||
		(x == 430 && y == 520) || (x == 481 && y == 7'd450) || (x == 7'd238 && y == 7'd353) ||
		(x == 7'd35 && y == 298) || (x == 7'd297 && y == 7'd622) || (x == 7'd439 && y == 7'd637) ||
		(x == 7'd501 && y == 529) || (x == 7'd292 && y == 227) || (x == 289 && y == 7'd111) ||
		(x == 7'd639 && y == 7'd49) || (x == 434 && y == 468) || (x == 38 && y == 7'd204) ||
		(x == 7'd579 && y == 7'd539) || (x == 7'd347 && y == 7'd461) || (x == 182 && y == 251) ||
		(x == 7'd214 && y == 7'd363) || (x == 7'd287 && y == 351) || (x == 321 && y == 387) ||
		(x == 7'd543 && y == 386) || (x == 68 && y == 70) || (x == 292 && y == 7'd617) ||
		(x == 7'd519 && y == 7'd286) || (x == 7'd132 && y == 428) || (x == 554 && y == 350) ||
		(x == 409 && y == 7'd283) || (x == 7'd572 && y == 269) || (x == 7'd330 && y == 7'd514) ||
		(x == 7'd418 && y == 7'd271) || (x == 7'd511 && y == 395) || (x == 7'd145 && y == 165) ||
		(x == 7'd167 && y == 7'd396) || (x == 7'd170 && y == 7'd298) || (x == 7'd251 && y == 382) ||
		(x == 568 && y == 272) || (x == 7'd376 && y == 297) || (x == 7'd450 && y == 436) ||
		(x == 7'd286 && y == 532) || (x == 7'd286 && y == 494) || (x == 7'd172 && y == 73) ||
		(x == 7'd136 && y == 119) || (x == 341 && y == 7'd537) || (x == 7'd624 && y == 7'd583) ||
		(x == 7'd164 && y == 229) || (x == 7'd285 && y == 7'd195) || (x == 7'd303 && y == 7'd253) ||
		(x == 146 && y == 7'd509) || (x == 197 && y == 222) || (x == 181 && y == 630) ||
		(x == 7'd498 && y == 7'd184) || (x == 195 && y == 7'd595) || (x == 629 && y == 7'd300) ||
		(x == 13 && y == 7'd116) || (x == 170 && y == 7'd268) || (x == 7'd160 && y == 7'd470) ||
		(x == 142 && y == 429) || (x == 7'd230 && y == 458) || (x == 322 && y == 7'd592) ||
		(x == 221 && y == 7'd344) || (x == 516 && y == 511) || (x == 7'd281 && y == 404) ||
		(x == 7'd509 && y == 506) || (x == 7'd227 && y == 147) || (x == 7'd444 && y == 7'd512) ||
		(x == 542 && y == 7'd514) || (x == 208 && y == 7'd476) || (x == 7'd569 && y == 383) ||
		(x == 571 && y == 220) || (x == 181 && y == 475) || (x == 7'd300 && y == 7'd158) ||
		(x == 451 && y == 597) || (x == 283 && y == 7'd498) || (x == 7'd122 && y == 7'd466) ||
		(x == 7'd534 && y == 7'd126) || (x == 639 && y == 307) || (x == 7'd465 && y == 7'd510) ||
		(x == 193 && y == 7'd607) || (x == 7'd370 && y == 304) || (x == 7'd399 && y == 195) ||
		(x == 329 && y == 7'd378) || (x == 255 && y == 7'd310) || (x == 266 && y == 7'd106) ||
		(x == 7'd215 && y == 303) || (x == 7'd440 && y == 7'd146) || (x == 499 && y == 7'd568) ||
		(x == 7'd535 && y == 329) || (x == 286 && y == 400) || (x == 7'd192 && y == 7'd198) ||
		(x == 7'd174 && y == 557) || (x == 321 && y == 332) || (x == 7'd90 && y == 453) ||
		(x == 7'd634 && y == 7'd490) || (x == 165 && y == 7'd424) || (x == 129 && y == 7'd526) ||
		(x == 317 && y == 7'd439) || (x == 7'd634 && y == 7'd194) || (x == 82 && y == 7'd595) ||
		(x == 179 && y == 7'd592) || (x == 267 && y == 467) || (x == 528 && y == 638) ||
		(x == 7'd407 && y == 7'd379) || (x == 562 && y == 618) || (x == 372 && y == 370) ||
		(x == 444 && y == 7'd612) || (x == 7'd242 && y == 7'd476) || (x == 7'd175 && y == 511) ||
		(x == 7'd377 && y == 7'd468) || (x == 446 && y == 151) || (x == 615 && y == 545) ||
		(x == 7'd565 && y == 568) || (x == 318 && y == 7'd244) || (x == 404 && y == 204) ||
		(x == 7'd527 && y == 7'd315) || (x == 7'd109 && y == 49) || (x == 7'd425 && y == 7'd468) ||
		(x == 496 && y == 503) || (x == 503 && y == 7'd316) || (x == 7'd622 && y == 7'd244) ||
		(x == 7'd373 && y == 198) || (x == 165 && y == 7'd173) || (x == 414 && y == 7'd9) ||
		(x == 7'd43 && y == 7'd261) || (x == 7'd178 && y == 7'd423) || (x == 249 && y == 441) ||
		(x == 7'd369 && y == 7'd261) || (x == 7'd322 && y == 392) || (x == 7'd227 && y == 7'd619) ||
		(x == 7'd265 && y == 7'd169) || (x == 208 && y == 7'd88) || (x == 7'd123 && y == 466) ||
		(x == 463 && y == 7'd121) || (x == 221 && y == 533) || (x == 21 && y == 7'd132) ||
		(x == 551 && y == 262) || (x == 70 && y == 7'd419) || (x == 7'd215 && y == 591) ||
		(x == 7'd607 && y == 7'd367) || (x == 7'd403 && y == 233) || (x == 73 && y == 7'd588) ||
		(x == 593 && y == 7'd581) || (x == 7'd342 && y == 384) || (x == 7'd532 && y == 7'd545) ||
		(x == 7'd521 && y == 7'd577) || (x == 492 && y == 7'd640) || (x == 7'd305 && y == 7'd513) ||
		(x == 7'd424 && y == 114) || (x == 283 && y == 392) || (x == 529 && y == 7'd219) ||
		(x == 192 && y == 7'd72) || (x == 7'd579 && y == 373) || (x == 7'd289 && y == 39) ||
		(x == 310 && y == 7'd249) || (x == 7'd474 && y == 7'd460) || (x == 7'd537 && y == 7'd263) ||
		(x == 501 && y == 7'd486) || (x == 235 && y == 7'd411) || (x == 7'd135 && y == 230) ||
		(x == 7'd444 && y == 7'd12) || (x == 7'd579 && y == 7'd186) || (x == 612 && y == 551) ||
		(x == 469 && y == 7'd206) || (x == 248 && y == 7'd172) || (x == 7'd560 && y == 445) ||
		(x == 7'd627 && y == 7'd634) || (x == 602 && y == 7'd143) || (x == 199 && y == 7'd395) ||
		(x == 204 && y == 7'd319) || (x == 364 && y == 7'd379) || (x == 7'd262 && y == 7'd493) ||
		(x == 517 && y == 460) || (x == 530 && y == 7'd634) || (x == 7'd54 && y == 205) ||
		(x == 37 && y == 7'd14) || (x == 7'd155 && y == 7'd258) || (x == 15 && y == 7'd276) ||
		(x == 319 && y == 7'd132) || (x == 401 && y == 131) || (x == 7'd429 && y == 581) ||
		(x == 7'd475 && y == 233) || (x == 7'd484 && y == 7'd400) || (x == 156 && y == 7'd442) ||
		(x == 458 && y == 159) || (x == 7'd569 && y == 429) || (x == 505 && y == 7'd582) ||
		(x == 7'd621 && y == 120) || (x == 7'd84 && y == 7'd507) || (x == 7'd133 && y == 430) ||
		(x == 7'd322 && y == 383) || (x == 7'd581 && y == 58) || (x == 564 && y == 347) ||
		(x == 7'd2 && y == 303) || (x == 198 && y == 7'd557) || (x == 7'd141 && y == 7'd335) ||
		(x == 7'd195 && y == 7'd434) || (x == 470 && y == 7'd173) || (x == 161 && y == 7'd494) ||
		(x == 292 && y == 339) || (x == 7'd220 && y == 7'd412) || (x == 596 && y == 215) ||
		(x == 7'd197 && y == 421) || (x == 599 && y == 246) || (x == 274 && y == 7'd374) ||
		(x == 620 && y == 222) || (x == 7'd451 && y == 7'd162) || (x == 245 && y == 7'd534) ||
		(x == 454 && y == 243) || (x == 418 && y == 7'd79) || (x == 7'd211 && y == 539) ||
		(x == 70 && y == 7'd548) || (x == 7'd263 && y == 7'd405) || (x == 7'd62 && y == 375) ||
		(x == 70 && y == 7'd363) || (x == 7'd171 && y == 275) || (x == 7'd600 && y == 624) ||
		(x == 7'd421 && y == 7'd385) || (x == 178 && y == 7'd544) || (x == 7'd78 && y == 194) ||
		(x == 287 && y == 7'd39) || (x == 242 && y == 293) || (x == 387 && y == 7'd457) ||
		(x == 383 && y == 7'd53) || (x == 7'd252 && y == 7'd282) || (x == 245 && y == 553) ||
		(x == 7'd526 && y == 7'd370) || (x == 159 && y == 410) || (x == 7'd355 && y == 189) ||
		(x == 601 && y == 583) || (x == 407 && y == 279) || (x == 7'd283 && y == 7'd269) ||
		(x == 398 && y == 7'd498) || (x == 389 && y == 7'd205) || (x == 137 && y == 534) ||
		(x == 77 && y == 7'd235) || (x == 7'd265 && y == 504) || (x == 7'd66 && y == 7'd477) ||
		(x == 187 && y == 7'd472) || (x == 7'd148 && y == 7'd632) || (x == 616 && y == 7'd182) ||
		(x == 7'd56 && y == 442) || (x == 7'd430 && y == 7'd254) || (x == 7'd17 && y == 7'd373) ||
		(x == 215 && y == 314) || (x == 7'd628 && y == 7'd622) || (x == 258 && y == 7'd474) ||
		(x == 99 && y == 7'd304) || (x == 468 && y == 7'd84) || (x == 534 && y == 7'd102) ||
		(x == 7'd392 && y == 575) || (x == 605 && y == 546) || (x == 7'd475 && y == 616) ||
		(x == 7'd130 && y == 7'd484) || (x == 7'd104 && y == 7'd353) || (x == 7'd271 && y == 34) ||
		(x == 7'd318 && y == 235) || (x == 48 && y == 7'd609) || (x == 383 && y == 149) ||
		(x == 270 && y == 351) || (x == 7'd261 && y == 7'd325) || (x == 7'd389 && y == 7'd153) ||
		(x == 7'd345 && y == 7'd403) || (x == 7'd413 && y == 7'd173) || (x == 543 && y == 367) ||
		(x == 7'd214 && y == 7'd95) || (x == 7'd565 && y == 7'd384) || (x == 549 && y == 7'd588) ||
		(x == 7'd400 && y == 504) || (x == 7'd342 && y == 7'd600) || (x == 7'd188 && y == 7'd634) ||
		(x == 221 && y == 7'd119) || (x == 7'd269 && y == 541) || (x == 614 && y == 7'd452) ||
		(x == 7'd223 && y == 7'd545) || (x == 7'd375 && y == 7'd493) || (x == 7'd190 && y == 7'd356) ||
		(x == 7'd611 && y == 7'd427) || (x == 7'd626 && y == 7'd249) || (x == 7'd372 && y == 85) ||
		(x == 7'd270 && y == 7'd239) || (x == 7'd370 && y == 479) || (x == 413 && y == 317) ||
		(x == 7'd554 && y == 95) || (x == 7'd485 && y == 7'd405) || (x == 7'd187 && y == 7'd379) ||
		(x == 553 && y == 478) || (x == 7'd338 && y == 7'd444) || (x == 7'd451 && y == 544) ||
		(x == 7'd60 && y == 570) || (x == 191 && y == 292) || (x == 545 && y == 7'd281) ||
		(x == 614 && y == 7'd484) || (x == 7'd476 && y == 7'd272) || (x == 373 && y == 7'd146) ||
		(x == 7'd269 && y == 155) || (x == 215 && y == 7'd337) || (x == 260 && y == 7'd529) ||
		(x == 7'd636 && y == 7'd147) || (x == 129 && y == 7'd168) || (x == 631 && y == 7'd456) ||
		(x == 410 && y == 216) || (x == 239 && y == 149) || (x == 7'd150 && y == 7'd260) ||
		(x == 559 && y == 7'd22) || (x == 7'd376 && y == 428) || (x == 7'd132 && y == 7'd134) ||
		(x == 64 && y == 7'd376) || (x == 7'd541 && y == 7'd381) || (x == 537 && y == 7'd555) ||
		(x == 314 && y == 228) || (x == 7'd466 && y == 153) || (x == 396 && y == 7'd326) ||
		(x == 395 && y == 296) || (x == 7'd516 && y == 7'd252) || (x == 7'd186 && y == 7'd623) ||
		(x == 7'd111 && y == 7'd159) || (x == 619 && y == 7'd9) || (x == 421 && y == 7'd165) ||
		(x == 7'd54 && y == 7'd40) || (x == 7'd5 && y == 7'd503) || (x == 7'd473 && y == 7'd401) ||
		(x == 7'd9 && y == 24) || (x == 600 && y == 321) || (x == 530 && y == 496) ||
		(x == 7'd85 && y == 543) || (x == 7'd72 && y == 7'd411) || (x == 213 && y == 7'd415) ||
		(x == 549 && y == 7'd184) || (x == 7'd608 && y == 7'd35) || (x == 7'd51 && y == 347) ||
		(x == 298 && y == 595) || (x == 199 && y == 502) || (x == 139 && y == 7'd81) ||
		(x == 7'd503 && y == 7'd168) || (x == 7'd348 && y == 7'd366) || (x == 7'd492 && y == 441) ||
		(x == 7'd376 && y == 7'd167) || (x == 7'd434 && y == 7'd516) || (x == 7'd502 && y == 7'd330) ||
		(x == 7'd524 && y == 169) || (x == 7'd138 && y == 7'd142) || (x == 7'd146 && y == 7'd506) ||
		(x == 7'd140 && y == 7'd469) || (x == 67 && y == 105) || (x == 7'd80 && y == 405) ||
		(x == 293 && y == 7'd336) || (x == 505 && y == 567) || (x == 446 && y == 599) ||
		(x == 7'd11 && y == 7'd345) || (x == 278 && y == 558) || (x == 7'd599 && y == 7'd344) ||
		(x == 189 && y == 7'd220) || (x == 7'd347 && y == 121) || (x == 273 && y == 7'd575) ||
		(x == 7'd535 && y == 163) || (x == 136 && y == 403) || (x == 112 && y == 7'd373) ||
		(x == 7'd345 && y == 7'd338) || (x == 7'd147 && y == 7'd269) || (x == 7'd82 && y == 354) ||
		(x == 7'd633 && y == 7'd209) || (x == 308 && y == 7'd23) || (x == 591 && y == 7'd593) ||
		(x == 7'd306 && y == 493) || (x == 593 && y == 7'd408) || (x == 7'd151 && y == 7'd139) ||
		(x == 76 && y == 7'd435) || (x == 7'd297 && y == 7'd435) || (x == 7'd526 && y == 7'd208) ||
		(x == 350 && y == 213) || (x == 7'd408 && y == 122) || (x == 7'd516 && y == 7'd289) ||
		(x == 432 && y == 7'd596) || (x == 7'd455 && y == 7'd368) || (x == 564 && y == 7'd46) ||
		(x == 221 && y == 372) || (x == 7'd442 && y == 19) || (x == 318 && y == 7'd56) ||
		(x == 7'd287 && y == 7'd468) || (x == 347 && y == 7'd557) || (x == 237 && y == 208) ||
		(x == 7'd12 && y == 392) || (x == 7'd608 && y == 129) || (x == 7'd425 && y == 169) ||
		(x == 304 && y == 187) || (x == 7'd499 && y == 108) || (x == 148 && y == 472) ||
		(x == 526 && y == 7'd550) || (x == 100 && y == 7'd361) || (x == 7'd619 && y == 7'd478) ||
		(x == 413 && y == 566) || (x == 7'd203 && y == 7'd272) || (x == 158 && y == 475) ||
		(x == 7'd377 && y == 435) || (x == 7'd254 && y == 7'd377) || (x == 7'd194 && y == 7'd368) ||
		(x == 516 && y == 326) || (x == 7'd176 && y == 7'd525) || (x == 7'd609 && y == 7'd7) ||
		(x == 331 && y == 580) || (x == 65 && y == 7'd296) || (x == 137 && y == 259) ||
		(x == 186 && y == 7'd99) || (x == 7'd188 && y == 204) || (x == 605 && y == 527) ||
		(x == 549 && y == 7'd26) || (x == 341 && y == 315) || (x == 7'd448 && y == 7'd630) ||
		(x == 7'd402 && y == 221) || (x == 7'd172 && y == 558) || (x == 7'd162 && y == 7'd248) ||
		(x == 311 && y == 7'd281) || (x == 409 && y == 619) || (x == 7'd304 && y == 7'd354) ||
		(x == 7'd555 && y == 7'd633) || (x == 7'd530 && y == 46) || (x == 157 && y == 543) ||
		(x == 512 && y == 553) || (x == 219 && y == 599) || (x == 524 && y == 7'd458) ||
		(x == 134 && y == 559) || (x == 390 && y == 7'd226) || (x == 7'd571 && y == 7'd85) ||
		(x == 7'd268 && y == 7'd149) || (x == 577 && y == 7'd237) || (x == 7'd114 && y == 7'd400) ||
		(x == 7'd404 && y == 183) || (x == 7'd328 && y == 7'd396) || (x == 7'd199 && y == 7'd526) ||
		(x == 7'd101 && y == 563) || (x == 423 && y == 228) || (x == 7'd575 && y == 278) ||
		(x == 7'd380 && y == 7'd257) || (x == 7'd536 && y == 7'd158) || (x == 244 && y == 210) ||
		(x == 566 && y == 297) || (x == 7'd530 && y == 7'd309) || (x == 104 && y == 7'd515) ||
		(x == 7'd134 && y == 7'd586) || (x == 517 && y == 485) || (x == 7'd457 && y == 192) ||
		(x == 7'd382 && y == 105) || (x == 7'd456 && y == 7'd512) || (x == 7'd532 && y == 220) ||
		(x == 132 && y == 7'd323) || (x == 7'd9 && y == 129) || (x == 7'd387 && y == 7'd222) ||
		(x == 7'd127 && y == 260) || (x == 338 && y == 511) || (x == 223 && y == 290) ||
		(x == 7'd212 && y == 7'd247) || (x == 7'd526 && y == 7'd549) || (x == 380 && y == 315) ||
		(x == 394 && y == 7'd200) || (x == 534 && y == 175) || (x == 606 && y == 578) ||
		(x == 7'd454 && y == 513) || (x == 511 && y == 155) || (x == 7'd152 && y == 7'd393) ||
		(x == 186 && y == 295) || (x == 136 && y == 7'd216) || (x == 469 && y == 7'd620) ||
		(x == 7'd190 && y == 107) || (x == 7'd393 && y == 75) || (x == 7'd105 && y == 7'd300) ||
		(x == 7'd386 && y == 7'd454) || (x == 421 && y == 388) || (x == 402 && y == 586) ||
		(x == 638 && y == 7'd482) || (x == 7'd14 && y == 7'd61) || (x == 7'd166 && y == 7'd100) ||
		(x == 7'd186 && y == 582) || (x == 7'd556 && y == 7'd510) || (x == 476 && y == 328) ||
		(x == 7'd55 && y == 207) || (x == 7'd623 && y == 7'd516) || (x == 261 && y == 632) ||
		(x == 320 && y == 7'd606) || (x == 7'd108 && y == 475) || (x == 256 && y == 168) ||
		(x == 7'd433 && y == 7'd131) || (x == 7'd136 && y == 7'd421) || (x == 218 && y == 7'd477) ||
		(x == 7'd547 && y == 7'd603) || (x == 328 && y == 462) || (x == 7'd524 && y == 7'd495) ||
		(x == 7'd358 && y == 7'd77) || (x == 370 && y == 7'd406) || (x == 7'd228 && y == 456) ||
		(x == 92 && y == 7'd113) || (x == 351 && y == 7'd633) || (x == 7'd365 && y == 7'd121) ||
		(x == 359 && y == 243) || (x == 7'd173 && y == 7'd228) || (x == 604 && y == 640) ||
		(x == 480 && y == 7'd151) || (x == 259 && y == 432) || (x == 535 && y == 7'd197) ||
		(x == 7'd66 && y == 316) || (x == 309 && y == 7'd435) || (x == 326 && y == 474) ||
		(x == 7'd518 && y == 586) || (x == 7'd638 && y == 7'd178) || (x == 360 && y == 616) ||
		(x == 7'd69 && y == 136) || (x == 7'd316 && y == 7'd13) || (x == 368 && y == 346) ||
		(x == 512 && y == 339) || (x == 576 && y == 7'd539) || (x == 318 && y == 7'd632) ||
		(x == 7'd122 && y == 577) || (x == 337 && y == 470) || (x == 227 && y == 358) ||
		(x == 137 && y == 7'd540) || (x == 169 && y == 183) || (x == 7'd246 && y == 7'd610) ||
		(x == 613 && y == 324) || (x == 194 && y == 281) || (x == 204 && y == 7'd613) ||
		(x == 7'd314 && y == 7'd198) || (x == 7'd282 && y == 217) || (x == 7'd293 && y == 477) ||
		(x == 536 && y == 7'd474) || (x == 7'd414 && y == 7'd466) || (x == 131 && y == 588) ||
		(x == 7'd504 && y == 441) || (x == 7'd395 && y == 7'd238) || (x == 7'd581 && y == 176) ||
		(x == 7'd410 && y == 294) || (x == 7'd463 && y == 344) || (x == 7'd520 && y == 7'd602) ||
		(x == 7'd426 && y == 7'd456) || (x == 186 && y == 7'd220) || (x == 215 && y == 7'd420) ||
		(x == 583 && y == 250) || (x == 594 && y == 397) || (x == 7'd325 && y == 7'd137) ||
		(x == 162 && y == 7'd162) || (x == 7'd81 && y == 7'd98) || (x == 7'd461 && y == 7'd305) ||
		(x == 7'd268 && y == 37) || (x == 7'd272 && y == 7'd568) || (x == 550 && y == 7'd360) ||
		(x == 7'd314 && y == 213) || (x == 7'd398 && y == 483) || (x == 89 && y == 7'd39) ||
		(x == 219 && y == 7'd583) || (x == 7'd496 && y == 7'd603) || (x == 7'd509 && y == 433) ||
		(x == 7'd461 && y == 350) || (x == 7'd212 && y == 7'd0) || (x == 355 && y == 7'd506) ||
		(x == 521 && y == 185) || (x == 7'd420 && y == 7'd529) || (x == 7'd373 && y == 7'd319) ||
		(x == 443 && y == 7'd551) || (x == 7'd218 && y == 198) || (x == 7'd299 && y == 627) ||
		(x == 7'd262 && y == 7'd285) || (x == 7'd506 && y == 7'd489) || (x == 7'd146 && y == 7'd196) ||
		(x == 7'd231 && y == 313) || (x == 7'd366 && y == 7'd20) || (x == 370 && y == 7'd377) ||
		(x == 499 && y == 424) || (x == 427 && y == 248) || (x == 7'd285 && y == 307) ||
		(x == 7'd249 && y == 239) || (x == 7'd482 && y == 7'd261) || (x == 7'd346 && y == 7'd481) ||
		(x == 343 && y == 173) || (x == 7'd631 && y == 7'd442) || (x == 7'd193 && y == 7'd174) ||
		(x == 7'd460 && y == 489) || (x == 7'd100 && y == 259) || (x == 134 && y == 375) ||
		(x == 256 && y == 7'd72) || (x == 7'd4 && y == 7'd482) || (x == 7'd135 && y == 7'd362) ||
		(x == 7'd634 && y == 366) || (x == 7'd486 && y == 7'd299) || (x == 638 && y == 7'd178) ||
		(x == 7'd382 && y == 7'd17) || (x == 170 && y == 7'd140) || (x == 538 && y == 7'd319) ||
		(x == 7'd94 && y == 175) || (x == 199 && y == 7'd252) || (x == 286 && y == 547) ||
		(x == 631 && y == 511) || (x == 420 && y == 273) || (x == 7'd259 && y == 231) ||
		(x == 7'd429 && y == 168) || (x == 7'd398 && y == 7'd23) || (x == 7'd609 && y == 492) ||
		(x == 7'd118 && y == 163) || (x == 355 && y == 7'd264) || (x == 7'd309 && y == 7'd105) ||
		(x == 291 && y == 7'd52) || (x == 199 && y == 7'd239) || (x == 7'd492 && y == 7'd513) ||
		(x == 390 && y == 617) || (x == 118 && y == 7'd290) || (x == 355 && y == 589) ||
		(x == 7'd227 && y == 7'd590) || (x == 7'd514 && y == 7'd202) || (x == 7'd176 && y == 7'd611) ||
		(x == 338 && y == 435) || (x == 516 && y == 250) || (x == 463 && y == 303) ||
		(x == 7'd135 && y == 607) || (x == 443 && y == 7'd488) || (x == 3 && y == 7'd195) ||
		(x == 265 && y == 7'd511) || (x == 7'd575 && y == 7'd554) || (x == 7'd183 && y == 629) ||
		(x == 595 && y == 7'd510) || (x == 7'd287 && y == 457) || (x == 7'd617 && y == 7'd256) ||
		(x == 230 && y == 259) || (x == 419 && y == 7'd357) || (x == 7'd595 && y == 7'd54) ||
		(x == 7'd370 && y == 7'd10) || (x == 7'd417 && y == 7'd502) || (x == 7'd235 && y == 557) ||
		(x == 7'd30 && y == 14) || (x == 145 && y == 398) || (x == 7'd324 && y == 7'd559) ||
		(x == 7'd534 && y == 7'd635) || (x == 7'd428 && y == 546) || (x == 7'd382 && y == 7'd245) ||
		(x == 570 && y == 7'd388) || (x == 398 && y == 7'd221) || (x == 348 && y == 577) ||
		(x == 7'd377 && y == 7'd267) || (x == 542 && y == 7'd147) || (x == 499 && y == 7'd358) ||
		(x == 552 && y == 393) || (x == 7'd527 && y == 7'd498) || (x == 7'd630 && y == 500) ||
		(x == 113 && y == 7'd12) || (x == 7'd252 && y == 7'd578) || (x == 7'd590 && y == 7'd299) ||
		(x == 7'd623 && y == 116) || (x == 156 && y == 460) || (x == 7'd89 && y == 183) ||
		(x == 529 && y == 200) || (x == 439 && y == 254) || (x == 7'd387 && y == 7'd156) ||
		(x == 445 && y == 7'd390) || (x == 97 && y == 7'd238) || (x == 7'd624 && y == 7'd119) ||
		(x == 479 && y == 7'd74) || (x == 357 && y == 7'd23) || (x == 590 && y == 7'd216) ||
		(x == 139 && y == 7'd51) || (x == 221 && y == 7'd458) || (x == 7'd519 && y == 7'd279) ||
		(x == 7'd301 && y == 553) || (x == 7'd225 && y == 485) || (x == 7'd321 && y == 7'd306) ||
		(x == 7'd269 && y == 7'd297) || (x == 7'd612 && y == 212) || (x == 7'd172 && y == 222) ||
		(x == 7'd431 && y == 619) || (x == 562 && y == 7'd281) || (x == 7'd501 && y == 579) ||
		(x == 329 && y == 7'd336) || (x == 102 && y == 7'd360) || (x == 7'd617 && y == 7'd558) ||
		(x == 340 && y == 7'd308) || (x == 332 && y == 7'd126) || (x == 420 && y == 377) ||
		(x == 7'd427 && y == 7'd85) || (x == 7'd617 && y == 7'd599) || (x == 7'd150 && y == 7'd175) ||
		(x == 377 && y == 277) || (x == 7'd520 && y == 7'd130) || (x == 217 && y == 417) ||
		(x == 7'd373 && y == 7'd352) || (x == 543 && y == 7'd513) || (x == 7'd216 && y == 7'd144) ||
		(x == 390 && y == 7'd546) || (x == 587 && y == 217) || (x == 7'd237 && y == 307) ||
		(x == 630 && y == 451) || (x == 261 && y == 466) || (x == 7'd634 && y == 7'd355) ||
		(x == 416 && y == 7'd26) || (x == 7'd380 && y == 7'd152) || (x == 512 && y == 322) ||
		(x == 591 && y == 575) || (x == 335 && y == 7'd569) || (x == 7'd254 && y == 7'd358) ||
		(x == 68 && y == 7'd35) || (x == 476 && y == 7'd292) || (x == 495 && y == 7'd119) ||
		(x == 589 && y == 630) || (x == 7'd463 && y == 7'd157) || (x == 316 && y == 223) ||
		(x == 7'd545 && y == 189) || (x == 605 && y == 7'd361) || (x == 427 && y == 251) ||
		(x == 7'd229 && y == 208) || (x == 396 && y == 433) || (x == 335 && y == 279) ||
		(x == 7'd553 && y == 7'd566) || (x == 110 && y == 7'd171) || (x == 7'd232 && y == 638) ||
		(x == 331 && y == 7'd162) || (x == 14 && y == 7'd548) || (x == 7'd363 && y == 7'd505) ||
		(x == 255 && y == 7'd430) || (x == 280 && y == 396) || (x == 498 && y == 7'd535) ||
		(x == 7'd80 && y == 7'd370) || (x == 7'd72 && y == 346) || (x == 364 && y == 421) ||
		(x == 7'd506 && y == 284) || (x == 7'd31 && y == 7'd258) || (x == 376 && y == 7'd216) ||
		(x == 7'd295 && y == 632) || (x == 7'd599 && y == 144) || (x == 7'd519 && y == 451) ||
		(x == 7'd36 && y == 224) || (x == 7'd51 && y == 598) || (x == 189 && y == 7'd170) ||
		(x == 485 && y == 150) || (x == 7'd47 && y == 7'd537) || (x == 7'd448 && y == 7'd140) ||
		(x == 230 && y == 241) || (x == 7'd626 && y == 7'd398) || (x == 365 && y == 7'd537) ||
		(x == 7'd109 && y == 7'd373) || (x == 7'd427 && y == 378) || (x == 7'd69 && y == 115) ||
		(x == 153 && y == 400) || (x == 7'd484 && y == 443) || (x == 121 && y == 7'd269) ||
		(x == 7'd624 && y == 7'd192) || (x == 364 && y == 7'd402) || (x == 608 && y == 347) ||
		(x == 333 && y == 188) || (x == 623 && y == 533) || (x == 7'd172 && y == 7'd506) ||
		(x == 227 && y == 202) || (x == 447 && y == 7'd306) || (x == 7'd281 && y == 7'd389) ||
		(x == 426 && y == 7'd554) || (x == 7 && y == 7'd576) || (x == 7'd401 && y == 7'd195) ||
		(x == 526 && y == 200) || (x == 189 && y == 489) || (x == 7'd71 && y == 465) ||
		(x == 384 && y == 632) || (x == 7'd68 && y == 7'd141) || (x == 183 && y == 7'd323) ||
		(x == 7'd374 && y == 191) || (x == 7'd349 && y == 7'd114) || (x == 7'd119 && y == 475) ||
		(x == 7'd170 && y == 151) || (x == 7'd269 && y == 7'd143) || (x == 7'd477 && y == 7'd625) ||
		(x == 284 && y == 7'd426) || (x == 7'd157 && y == 388) || (x == 471 && y == 7'd348) ||
		(x == 92 && y == 7'd289) || (x == 7'd282 && y == 587) || (x == 334 && y == 483) ||
		(x == 7'd449 && y == 7'd135) || (x == 625 && y == 371) || (x == 7'd288 && y == 290) ||
		(x == 7'd578 && y == 7'd73) || (x == 7'd298 && y == 241) || (x == 162 && y == 7'd177) ||
		(x == 7'd249 && y == 75) || (x == 7'd453 && y == 480) || (x == 7'd255 && y == 7'd306) ||
		(x == 7'd168 && y == 7'd328) || (x == 553 && y == 376) || (x == 7'd93 && y == 7'd396) ||
		(x == 472 && y == 7'd39) || (x == 284 && y == 259) || (x == 7'd628 && y == 7'd635) ||
		(x == 7'd352 && y == 7'd562) || (x == 147 && y == 7'd457) || (x == 138 && y == 7'd543) ||
		(x == 524 && y == 7'd258) || (x == 7'd454 && y == 7'd3) || (x == 7'd472 && y == 7'd529) ||
		(x == 385 && y == 7'd425) || (x == 308 && y == 176) || (x == 558 && y == 282) ||
		(x == 7'd263 && y == 7'd570) || (x == 7'd20 && y == 7'd179) || (x == 7'd67 && y == 7'd244) ||
		(x == 7'd557 && y == 7'd250) || (x == 7'd24 && y == 192) || (x == 7'd212 && y == 480) ||
		(x == 173 && y == 268) || (x == 7'd58 && y == 336) || (x == 7'd384 && y == 510) ||
		(x == 362 && y == 307) || (x == 221 && y == 453) || (x == 7'd420 && y == 7'd513) ||
		(x == 522 && y == 7'd429) || (x == 533 && y == 623) || (x == 7'd156 && y == 583) ||
		(x == 554 && y == 458) || (x == 138 && y == 7'd270) || (x == 322 && y == 7'd381) ||
		(x == 7'd349 && y == 7'd290) || (x == 338 && y == 315) || (x == 328 && y == 462) ||
		(x == 582 && y == 308) || (x == 528 && y == 190) || (x == 7'd34 && y == 130) ||
		(x == 7'd182 && y == 7'd574) || (x == 7'd581 && y == 7'd419) || (x == 132 && y == 462) ||
		(x == 7'd315 && y == 7'd0) || (x == 440 && y == 7'd502) || (x == 7'd459 && y == 162) ||
		(x == 7'd347 && y == 7'd140) || (x == 459 && y == 7'd262) || (x == 7'd377 && y == 7'd12) ||
		(x == 46 && y == 7'd262) || (x == 7'd255 && y == 621) || (x == 7'd379 && y == 7'd262) ||
		(x == 7'd515 && y == 7'd396) || (x == 467 && y == 7'd601) || (x == 207 && y == 265) ||
		(x == 7'd629 && y == 99) || (x == 7'd180 && y == 7'd388) || (x == 7'd508 && y == 564) ||
		(x == 238 && y == 7'd307) || (x == 7'd246 && y == 7'd495) || (x == 478 && y == 533) ||
		(x == 7'd561 && y == 559) || (x == 7'd110 && y == 270) || (x == 7'd625 && y == 7'd295) ||
		(x == 147 && y == 434) || (x == 570 && y == 7'd169) || (x == 530 && y == 7'd358) ||
		(x == 349 && y == 7'd179) || (x == 7'd128 && y == 201) || (x == 7'd314 && y == 7'd638) ||
		(x == 194 && y == 158) || (x == 7'd226 && y == 383) || (x == 7'd529 && y == 2) ||
		(x == 291 && y == 492) || (x == 7'd400 && y == 7'd145) || (x == 7'd35 && y == 7'd500) ||
		(x == 7'd70 && y == 7'd541) || (x == 7'd613 && y == 379) || (x == 7'd240 && y == 159) ||
		(x == 167 && y == 7'd336) || (x == 7'd521 && y == 582) || (x == 7'd289 && y == 7'd343) ||
		(x == 7'd292 && y == 597) || (x == 190 && y == 495) || (x == 7'd244 && y == 7'd38) ||
		(x == 547 && y == 7'd445) || (x == 338 && y == 547) || (x == 7'd360 && y == 7'd513) ||
		(x == 7'd339 && y == 238) || (x == 7'd538 && y == 7'd509) || (x == 590 && y == 7'd470) ||
		(x == 7'd74 && y == 305) || (x == 489 && y == 262) || (x == 7'd637 && y == 298) ||
		(x == 352 && y == 424) || (x == 535 && y == 510) || (x == 209 && y == 7'd292) ||
		(x == 7'd78 && y == 485) || (x == 334 && y == 7'd410) || (x == 7'd400 && y == 7'd450) ||
		(x == 256 && y == 616) || (x == 568 && y == 7'd181) || (x == 293 && y == 409) ||
		(x == 8 && y == 7'd572) || (x == 7'd562 && y == 445) || (x == 202 && y == 7'd161) ||
		(x == 577 && y == 450) || (x == 7'd278 && y == 7'd335) || (x == 277 && y == 390) ||
		(x == 7'd365 && y == 279) || (x == 7'd40 && y == 7'd502) || (x == 7'd192 && y == 7'd388) ||
		(x == 7'd13 && y == 7'd274) || (x == 598 && y == 7'd584) || (x == 7'd524 && y == 7'd575) ||
		(x == 7'd288 && y == 407) || (x == 7'd506 && y == 7'd284) || (x == 7'd556 && y == 620) ||
		(x == 7'd449 && y == 7'd229) || (x == 7'd242 && y == 161) || (x == 7'd393 && y == 295) ||
		(x == 338 && y == 216) || (x == 7'd583 && y == 7'd589) || (x == 7'd554 && y == 7'd341) ||
		(x == 7'd342 && y == 7'd424) || (x == 7'd310 && y == 270) || (x == 7'd494 && y == 3) ||
		(x == 7'd186 && y == 7'd471) || (x == 268 && y == 7'd123) || (x == 187 && y == 370) ||
		(x == 7'd633 && y == 7'd160) || (x == 7'd17 && y == 43) || (x == 313 && y == 7'd160) ||
		(x == 7'd165 && y == 7'd316) || (x == 7'd56 && y == 7'd369) || (x == 358 && y == 396) ||
		(x == 572 && y == 260) || (x == 495 && y == 599) || (x == 585 && y == 7'd557) ||
		(x == 7'd447 && y == 381) || (x == 567 && y == 7'd285) || (x == 251 && y == 7'd47) ||
		(x == 225 && y == 467) || (x == 7'd295 && y == 89) || (x == 7'd147 && y == 7'd432) ||
		(x == 204 && y == 7'd628) || (x == 7'd617 && y == 7'd628) || (x == 7'd236 && y == 419) ||
		(x == 7'd378 && y == 7'd575) || (x == 302 && y == 7'd280) || (x == 7'd456 && y == 126) ||
		(x == 322 && y == 591) || (x == 209 && y == 7'd18) || (x == 538 && y == 616) ||
		(x == 304 && y == 167) || (x == 7'd395 && y == 7'd512) || (x == 524 && y == 7'd25) ||
		(x == 7'd133 && y == 7'd521) || (x == 7'd14 && y == 7'd142) || (x == 286 && y == 253) ||
		(x == 7'd119 && y == 7'd316) || (x == 7'd93 && y == 7'd343) || (x == 7'd353 && y == 7'd303) ||
		(x == 50 && y == 7'd0) || (x == 7'd401 && y == 188) || (x == 180 && y == 7'd402) ||
		(x == 7'd348 && y == 7'd309) || (x == 384 && y == 7'd83) || (x == 7'd637 && y == 7'd84) ||
		(x == 7'd181 && y == 467) || (x == 87 && y == 7'd134) || (x == 474 && y == 7'd331) ||
		(x == 630 && y == 592) || (x == 119 && y == 7'd415) || (x == 7'd262 && y == 7'd303) ||
		(x == 7'd263 && y == 7'd420) || (x == 7'd79 && y == 7'd378) || (x == 7'd164 && y == 7'd373) ||
		(x == 444 && y == 445) || (x == 203 && y == 7'd152) || (x == 7'd623 && y == 448) ||
		(x == 7'd2 && y == 551) || (x == 156 && y == 7'd610) || (x == 466 && y == 7'd431) ||
		(x == 640 && y == 7'd466) || (x == 7'd291 && y == 7'd59) || (x == 7'd244 && y == 7'd94) ||
		(x == 468 && y == 150) || (x == 7'd283 && y == 7'd303) || (x == 475 && y == 7'd103) ||
		(x == 7'd212 && y == 361) || (x == 7'd351 && y == 345) || (x == 7'd586 && y == 7'd428) ||
		(x == 138 && y == 431) || (x == 535 && y == 451) || (x == 7'd128 && y == 347) ||
		(x == 144 && y == 527) || (x == 7'd274 && y == 226) || (x == 336 && y == 135) ||
		(x == 7'd378 && y == 257) || (x == 7'd453 && y == 156) || (x == 278 && y == 7'd625) ||
		(x == 210 && y == 7'd446) || (x == 7'd496 && y == 7'd449) || (x == 257 && y == 315) ||
		(x == 7'd514 && y == 7'd72) || (x == 7'd507 && y == 589) || (x == 7'd31 && y == 7'd578) ||
		(x == 421 && y == 7'd163) || (x == 614 && y == 7'd585) || (x == 171 && y == 7'd213) ||
		(x == 370 && y == 7'd182) || (x == 7'd267 && y == 7'd550) || (x == 7'd428 && y == 7'd62) ||
		(x == 504 && y == 7'd53) || (x == 7'd273 && y == 7'd310) || (x == 200 && y == 394) ||
		(x == 118 && y == 7'd362) || (x == 7'd332 && y == 7'd614) || (x == 7'd137 && y == 7'd128) ||
		(x == 7'd7 && y == 7'd630) || (x == 7'd370 && y == 7'd291) || (x == 7'd245 && y == 7'd543) ||
		(x == 492 && y == 568) || (x == 554 && y == 7'd514) || (x == 7'd473 && y == 620) ||
		(x == 581 && y == 361) || (x == 7'd130 && y == 313) || (x == 7'd139 && y == 7'd426) ||
		(x == 385 && y == 7'd350) || (x == 99 && y == 7'd209) || (x == 7'd469 && y == 7'd348) ||
		(x == 7'd570 && y == 418) || (x == 319 && y == 199) || (x == 7'd499 && y == 529) ||
		(x == 453 && y == 7'd289) || (x == 296 && y == 133) || (x == 266 && y == 7'd241) ||
		(x == 7'd598 && y == 471) || (x == 636 && y == 342) || (x == 527 && y == 474) ||
		(x == 436 && y == 184) || (x == 7'd482 && y == 7'd527) || (x == 527 && y == 7'd606) ||
		(x == 590 && y == 7'd179) || (x == 7'd505 && y == 7'd508) || (x == 7'd210 && y == 7'd576) ||
		(x == 7'd116 && y == 61) || (x == 7'd633 && y == 7'd319) || (x == 366 && y == 420) ||
		(x == 7'd316 && y == 116) || (x == 7'd254 && y == 7'd280) || (x == 7'd305 && y == 513) ||
		(x == 7'd193 && y == 7'd268) || (x == 310 && y == 7'd455) || (x == 605 && y == 239) ||
		(x == 7'd164 && y == 631) || (x == 165 && y == 138) || (x == 545 && y == 318) ||
		(x == 7'd528 && y == 7'd501) || (x == 7'd332 && y == 251) || (x == 7'd140 && y == 7'd89) ||
		(x == 7'd340 && y == 437) || (x == 7'd93 && y == 168) || (x == 7'd441 && y == 7'd196) ||
		(x == 294 && y == 582) || (x == 7'd217 && y == 7'd499) || (x == 51 && y == 7'd385) ||
		(x == 52 && y == 7'd436) || (x == 7'd498 && y == 315) || (x == 7'd622 && y == 7'd433) ||
		(x == 326 && y == 7'd14) || (x == 7'd244 && y == 7'd288) || (x == 7'd432 && y == 7'd135) ||
		(x == 179 && y == 7'd203) || (x == 7'd444 && y == 461) || (x == 7'd589 && y == 442) ||
		(x == 468 && y == 7'd461) || (x == 7'd509 && y == 7'd174) || (x == 274 && y == 361) ||
		(x == 7'd12 && y == 519) || (x == 7'd92 && y == 7'd522) || (x == 510 && y == 502) ||
		(x == 7'd219 && y == 7'd391) || (x == 436 && y == 308) || (x == 7'd383 && y == 7'd560) ||
		(x == 7'd583 && y == 7'd186) || (x == 134 && y == 130) || (x == 218 && y == 7'd459) ||
		(x == 7'd355 && y == 7'd520) || (x == 356 && y == 253) || (x == 207 && y == 7'd517) ||
		(x == 7'd507 && y == 7'd632) || (x == 7'd574 && y == 7'd505) || (x == 77 && y == 7'd455) ||
		(x == 7'd500 && y == 7'd347) || (x == 7'd590 && y == 50) || (x == 7'd284 && y == 225) ||
		(x == 359 && y == 7'd300) || (x == 7'd545 && y == 7'd377) || (x == 7'd305 && y == 274) ||
		(x == 7'd41 && y == 535) || (x == 184 && y == 437) || (x == 7'd183 && y == 7'd252) ||
		(x == 148 && y == 203) || (x == 7'd519 && y == 7'd251) || (x == 7'd505 && y == 169) ||
		(x == 332 && y == 322) || (x == 7'd98 && y == 258) || (x == 582 && y == 513) ||
		(x == 179 && y == 7'd257) || (x == 457 && y == 188) || (x == 7'd78 && y == 622) ||
		(x == 379 && y == 7'd526) || (x == 79 && y == 50) || (x == 7'd296 && y == 7'd599) ||
		(x == 577 && y == 7'd411) || (x == 392 && y == 7'd125) || (x == 7'd216 && y == 7'd504) ||
		(x == 7'd225 && y == 71) || (x == 7'd337 && y == 7'd28) || (x == 7'd355 && y == 7'd333) ||
		(x == 271 && y == 7'd611) || (x == 117 && y == 7'd382) || (x == 7'd349 && y == 294) ||
		(x == 7'd194 && y == 7'd188) || (x == 7'd338 && y == 157) || (x == 520 && y == 7'd357) ||
		(x == 40 && y == 7'd597) || (x == 7'd314 && y == 82) || (x == 152 && y == 7'd602) ||
		(x == 572 && y == 174) || (x == 445 && y == 7'd224) || (x == 258 && y == 7'd83) ||
		(x == 398 && y == 7'd185) || (x == 7'd247 && y == 132) || (x == 7'd280 && y == 575) ||
		(x == 7'd528 && y == 7'd580) || (x == 7'd360 && y == 7'd615) || (x == 7'd135 && y == 7'd233) ||
		(x == 7'd551 && y == 7'd216) || (x == 7'd264 && y == 7'd322) || (x == 7'd206 && y == 7'd175) ||
		(x == 551 && y == 514) || (x == 7'd407 && y == 7'd564) || (x == 7'd210 && y == 241) ||
		(x == 7'd330 && y == 218) || (x == 7'd516 && y == 7'd541) || (x == 7'd396 && y == 7'd513) ||
		(x == 453 && y == 247) || (x == 7'd467 && y == 7'd363) || (x == 231 && y == 7'd115) ||
		(x == 372 && y == 213) || (x == 7'd35 && y == 323) || (x == 266 && y == 7'd438) ||
		(x == 7'd253 && y == 4) || (x == 7'd565 && y == 7'd199) || (x == 373 && y == 7'd12) ||
		(x == 160 && y == 7'd303) || (x == 7'd418 && y == 528) || (x == 7'd273 && y == 7'd526) ||
		(x == 212 && y == 406) || (x == 7'd480 && y == 7'd180) || (x == 581 && y == 322) ||
		(x == 50 && y == 7'd37) || (x == 7'd492 && y == 88) || (x == 7'd579 && y == 7'd455) ||
		(x == 7'd244 && y == 7'd216) || (x == 631 && y == 7'd174) || (x == 7'd244 && y == 7'd367) ||
		(x == 7'd376 && y == 7'd516) || (x == 7'd201 && y == 7'd459) || (x == 7'd473 && y == 562) ||
		(x == 7'd606 && y == 150) || (x == 261 && y == 7'd617) || (x == 171 && y == 7'd47) ||
		(x == 264 && y == 442) || (x == 557 && y == 389) || (x == 7'd453 && y == 7'd336) ||
		(x == 429 && y == 459) || (x == 7'd44 && y == 461) || (x == 7'd277 && y == 7'd55) ||
		(x == 7'd474 && y == 7'd8) || (x == 7'd103 && y == 7'd157) || (x == 387 && y == 7'd512) ||
		(x == 7'd193 && y == 7'd30) || (x == 7'd103 && y == 7'd23) || (x == 7'd102 && y == 7'd486) ||
		(x == 273 && y == 7'd460) || (x == 7'd475 && y == 7'd429) || (x == 289 && y == 546) ||
		(x == 7'd390 && y == 7'd186) || (x == 288 && y == 427) || (x == 7'd292 && y == 7'd350) ||
		(x == 211 && y == 297) || (x == 68 && y == 7'd520) || (x == 7'd135 && y == 423) ||
		(x == 7'd326 && y == 7'd113) || (x == 7'd480 && y == 615) || (x == 203 && y == 201) ||
		(x == 7'd208 && y == 7'd385) || (x == 7'd322 && y == 7'd138) || (x == 7'd109 && y == 303) ||
		(x == 7'd473 && y == 7'd173) || (x == 7'd213 && y == 440) || (x == 7'd582 && y == 7'd12) ||
		(x == 7'd249 && y == 7'd610) || (x == 7'd574 && y == 7'd391) || (x == 7'd614 && y == 321) ||
		(x == 340 && y == 153) || (x == 7'd486 && y == 442) || (x == 156 && y == 7'd100) ||
		(x == 466 && y == 7'd134) || (x == 342 && y == 7'd631) || (x == 7'd84 && y == 284) ||
		(x == 547 && y == 627) || (x == 137 && y == 7'd525) || (x == 7'd243 && y == 7'd262) ||
		(x == 7'd96 && y == 528) || (x == 7'd8 && y == 7'd440) || (x == 7'd288 && y == 424) ||
		(x == 533 && y == 7'd57) || (x == 498 && y == 468) || (x == 7'd3 && y == 7'd227) ||
		(x == 7'd461 && y == 412) || (x == 485 && y == 608) || (x == 361 && y == 7'd145) ||
		(x == 407 && y == 7'd67) || (x == 7'd106 && y == 113) || (x == 7'd487 && y == 7'd465) ||
		(x == 7'd480 && y == 7'd618) || (x == 7'd109 && y == 7'd197) || (x == 7'd580 && y == 566) ||
		(x == 7'd286 && y == 170) || (x == 377 && y == 7'd29) || (x == 256 && y == 546) ||
		(x == 7'd130 && y == 7'd265) || (x == 215 && y == 7'd298) || (x == 7'd539 && y == 170) ||
		(x == 466 && y == 7'd403) || (x == 157 && y == 317) || (x == 350 && y == 7'd593) ||
		(x == 625 && y == 405) || (x == 187 && y == 7'd312) || (x == 549 && y == 567) ||
		(x == 7'd316 && y == 7'd83) || (x == 7'd376 && y == 284) || (x == 27 && y == 7'd136) ||
		(x == 7'd422 && y == 7'd248) || (x == 7'd258 && y == 7'd329) || (x == 591 && y == 7'd638) ||
		(x == 7'd459 && y == 7'd48) || (x == 7'd18 && y == 7'd45) || (x == 7'd455 && y == 479) ||
		(x == 7'd352 && y == 535) || (x == 7'd516 && y == 7'd154) || (x == 7'd552 && y == 583) ||
		(x == 103 && y == 7'd229) || (x == 287 && y == 7'd557) || (x == 7'd574 && y == 115) ||
		(x == 7'd321 && y == 7'd581) || (x == 178 && y == 299) || (x == 474 && y == 7'd108) ||
		(x == 431 && y == 220) || (x == 7'd192 && y == 7'd137) || (x == 105 && y == 7'd356) ||
		(x == 364 && y == 314) || (x == 516 && y == 7'd608) || (x == 7'd417 && y == 214) ||
		(x == 7'd345 && y == 405) || (x == 436 && y == 386) || (x == 569 && y == 7'd413) ||
		(x == 338 && y == 197) || (x == 7'd106 && y == 7'd84) || (x == 375 && y == 7'd230) ||
		(x == 218 && y == 7'd186) || (x == 7'd190 && y == 181) || (x == 7'd65 && y == 7'd187) ||
		(x == 7'd628 && y == 334) || (x == 313 && y == 7'd81) || (x == 14 && y == 7'd210) ||
		(x == 369 && y == 7'd108) || (x == 469 && y == 7'd188) || (x == 199 && y == 565) ||
		(x == 281 && y == 7'd377) || (x == 318 && y == 7'd314) || (x == 7'd554 && y == 276) ||
		(x == 7'd514 && y == 7'd253) || (x == 7'd18 && y == 7'd281) || (x == 7'd295 && y == 7'd343) ||
		(x == 7'd577 && y == 7'd136) || (x == 7'd381 && y == 7'd284) || (x == 7'd350 && y == 111) ||
		(x == 7'd162 && y == 98) || (x == 7'd364 && y == 7'd601) || (x == 304 && y == 7'd293) ||
		(x == 419 && y == 7'd493) || (x == 530 && y == 371) || (x == 553 && y == 143) ||
		(x == 7'd152 && y == 7'd389) || (x == 495 && y == 600) || (x == 313 && y == 296) ||
		(x == 7'd200 && y == 7'd441) || (x == 347 && y == 7'd557) || (x == 334 && y == 498) ||
		(x == 174 && y == 7'd346) || (x == 187 && y == 450) || (x == 7'd496 && y == 7'd292) ||
		(x == 7'd369 && y == 388) || (x == 7'd332 && y == 7'd401) || (x == 7'd61 && y == 257) ||
		(x == 443 && y == 7'd110) || (x == 7'd360 && y == 125) || (x == 229 && y == 329) ||
		(x == 194 && y == 7'd506) || (x == 138 && y == 7'd43) || (x == 570 && y == 617) ||
		(x == 7'd365 && y == 7'd39) || (x == 452 && y == 7'd64) || (x == 7'd238 && y == 7'd402) ||
		(x == 7'd446 && y == 7'd388) || (x == 7'd547 && y == 7'd483) || (x == 469 && y == 7'd513) ||
		(x == 7'd67 && y == 396) || (x == 7'd482 && y == 387) || (x == 186 && y == 7'd601) ||
		(x == 292 && y == 7'd525) || (x == 515 && y == 7'd637) || (x == 7'd633 && y == 434) ||
		(x == 7'd365 && y == 7'd531) || (x == 7'd554 && y == 7'd249) || (x == 7'd467 && y == 378) ||
		(x == 419 && y == 275) || (x == 7'd375 && y == 7'd315) || (x == 249 && y == 7'd342) ||
		(x == 323 && y == 7'd247) || (x == 7'd326 && y == 7'd461) || (x == 7'd555 && y == 7'd226) ||
		(x == 7'd24 && y == 638) || (x == 209 && y == 231) || (x == 330 && y == 7'd377) ||
		(x == 231 && y == 7'd626) || (x == 570 && y == 141) || (x == 7'd523 && y == 323) ||
		(x == 7'd400 && y == 7'd627) || (x == 195 && y == 7'd70) || (x == 7'd458 && y == 7'd177) ||
		(x == 7'd292 && y == 7'd604) || (x == 7'd248 && y == 79) || (x == 7'd525 && y == 375) ||
		(x == 7'd342 && y == 86) || (x == 7'd324 && y == 7'd27) || (x == 109 && y == 7'd277) ||
		(x == 7'd327 && y == 7'd395) || (x == 7'd19 && y == 7'd558) || (x == 570 && y == 7'd53) ||
		(x == 568 && y == 7'd177) || (x == 7'd101 && y == 7'd258) || (x == 486 && y == 187) ||
		(x == 223 && y == 7'd338) || (x == 282 && y == 209) || (x == 7'd425 && y == 7'd355) ||
		(x == 163 && y == 7'd463) || (x == 7'd359 && y == 115) || (x == 562 && y == 224) ||
		(x == 623 && y == 7'd47) || (x == 69 && y == 7'd458) || (x == 7'd629 && y == 628) ||
		(x == 7'd16 && y == 62) || (x == 7'd310 && y == 545) || (x == 7'd330 && y == 638) ||
		(x == 174 && y == 7'd509) || (x == 7'd331 && y == 7'd216) || (x == 132 && y == 435) ||
		(x == 317 && y == 366) || (x == 7'd439 && y == 7'd17) || (x == 535 && y == 252) ||
		(x == 7'd448 && y == 293) || (x == 7'd323 && y == 7'd92) || (x == 291 && y == 7'd523) ||
		(x == 81 && y == 75) || (x == 225 && y == 7'd269) || (x == 625 && y == 7'd347) ||
		(x == 355 && y == 7'd248) || (x == 159 && y == 7'd540) || (x == 7'd444 && y == 7'd313) ||
		(x == 452 && y == 131) || (x == 225 && y == 7'd92) || (x == 7'd538 && y == 283) ||
		(x == 340 && y == 7'd541) || (x == 485 && y == 271) || (x == 7'd63 && y == 438) ||
		(x == 7'd496 && y == 7'd141) || (x == 639 && y == 7'd576) || (x == 163 && y == 241) ||
		(x == 548 && y == 7'd380) || (x == 381 && y == 285) || (x == 7'd138 && y == 42) ||
		(x == 7'd379 && y == 7'd451) || (x == 262 && y == 7'd84) || (x == 5 && y == 7'd224) ||
		(x == 7'd301 && y == 433) || (x == 7'd635 && y == 7'd38) || (x == 575 && y == 7'd148) ||
		(x == 309 && y == 224) || (x == 313 && y == 357) || (x == 7'd297 && y == 7'd623) ||
		(x == 7'd390 && y == 7'd394) || (x == 433 && y == 258) || (x == 420 && y == 7'd502) ||
		(x == 7'd243 && y == 7'd392) || (x == 7'd453 && y == 7'd517) || (x == 7'd12 && y == 500) ||
		(x == 7'd171 && y == 369) || (x == 7'd304 && y == 7'd395) || (x == 7'd159 && y == 473) ||
		(x == 7'd152 && y == 619) || (x == 7'd13 && y == 7'd551) || (x == 7'd47 && y == 7'd259) ||
		(x == 7'd534 && y == 7'd508) || (x == 7'd85 && y == 178) || (x == 527 && y == 245) ||
		(x == 7'd634 && y == 7'd438) || (x == 7'd478 && y == 607) || (x == 589 && y == 631) ||
		(x == 548 && y == 310) || (x == 7'd639 && y == 7'd81) || (x == 533 && y == 378) ||
		(x == 7'd175 && y == 406) || (x == 281 && y == 211) || (x == 7'd462 && y == 7'd45) ||
		(x == 7'd189 && y == 177) || (x == 7'd411 && y == 572) || (x == 7'd438 && y == 373) ||
		(x == 88 && y == 71) || (x == 7'd184 && y == 7'd528) || (x == 502 && y == 7'd94) ||
		(x == 200 && y == 7'd271) || (x == 134 && y == 7'd98) || (x == 540 && y == 537) ||
		(x == 442 && y == 7'd380) || (x == 7'd388 && y == 97) || (x == 7'd171 && y == 581) ||
		(x == 129 && y == 7'd320) || (x == 7'd21 && y == 521) || (x == 329 && y == 7'd17) ||
		(x == 7'd56 && y == 7'd506) || (x == 496 && y == 7'd316) || (x == 7'd550 && y == 7'd472) ||
		(x == 350 && y == 553) || (x == 7'd505 && y == 7'd64) || (x == 595 && y == 525) ||
		(x == 7'd402 && y == 7'd300) || (x == 531 && y == 577) || (x == 82 && y == 7'd111) ||
		(x == 7'd369 && y == 7'd565) || (x == 7'd239 && y == 236) || (x == 199 && y == 7'd311) ||
		(x == 7'd125 && y == 16) || (x == 7'd458 && y == 7'd43) || (x == 7'd526 && y == 7'd43) ||
		(x == 7'd237 && y == 7'd180) || (x == 7'd373 && y == 7'd317) || (x == 187 && y == 7'd125) ||
		(x == 338 && y == 593) || (x == 7'd6 && y == 7'd585) || (x == 278 && y == 413) ||
		(x == 7'd392 && y == 175) || (x == 7'd473 && y == 7'd553) || (x == 430 && y == 538) ||
		(x == 7'd590 && y == 7'd590) || (x == 7'd419 && y == 7'd499) || (x == 7'd159 && y == 7'd617) ||
		(x == 158 && y == 7'd204) || (x == 7'd449 && y == 274) || (x == 570 && y == 318) ||
		(x == 7'd502 && y == 542) || (x == 7'd17 && y == 65) || (x == 322 && y == 373) ||
		(x == 387 && y == 7'd512) || (x == 7'd521 && y == 7'd451) || (x == 529 && y == 7'd197) ||
		(x == 233 && y == 361) || (x == 7'd155 && y == 7'd395) || (x == 7'd40 && y == 319) ||
		(x == 313 && y == 7'd585) || (x == 204 && y == 7'd572) || (x == 580 && y == 7'd565) ||
		(x == 7'd558 && y == 7'd165) || (x == 398 && y == 269) || (x == 565 && y == 481) ||
		(x == 7'd316 && y == 7'd629) || (x == 7'd242 && y == 591) || (x == 543 && y == 382) ||
		(x == 338 && y == 7'd304) || (x == 7'd321 && y == 7'd446) || (x == 7'd319 && y == 460) ||
		(x == 90 && y == 7'd551) || (x == 540 && y == 479) || (x == 7'd623 && y == 7'd243) ||
		(x == 7'd500 && y == 7'd520) || (x == 364 && y == 565) || (x == 7'd406 && y == 7'd302) ||
		(x == 7'd184 && y == 7'd623) || (x == 359 && y == 7'd468) || (x == 7'd304 && y == 212) ||
		(x == 7'd472 && y == 7'd246) || (x == 268 && y == 335) || (x == 7'd328 && y == 277) ||
		(x == 7'd92 && y == 439) || (x == 634 && y == 185) || (x == 7'd322 && y == 7'd602) ||
		(x == 7'd514 && y == 382) || (x == 622 && y == 7'd18) || (x == 7'd276 && y == 7'd208) ||
		(x == 210 && y == 368) || (x == 292 && y == 7'd236) || (x == 7'd320 && y == 7'd266) ||
		(x == 287 && y == 514) || (x == 7'd467 && y == 291) || (x == 425 && y == 556) ||
		(x == 58 && y == 7'd124) || (x == 7'd425 && y == 441) || (x == 7'd502 && y == 7'd460) ||
		(x == 7'd345 && y == 7'd269) || (x == 7'd331 && y == 478) || (x == 34 && y == 7'd18) ||
		(x == 7'd317 && y == 273) || (x == 181 && y == 7'd297) || (x == 90 && y == 7'd141) ||
		(x == 7'd100 && y == 483) || (x == 637 && y == 570) || (x == 469 && y == 490) ||
		(x == 53 && y == 27) || (x == 205 && y == 361) || (x == 559 && y == 161) ||
		(x == 484 && y == 7'd597) || (x == 156 && y == 7'd133) || (x == 552 && y == 7'd8) ||
		(x == 7'd383 && y == 7'd20) || (x == 7'd313 && y == 7'd530) || (x == 7'd318 && y == 589) ||
		(x == 7'd259 && y == 586) || (x == 264 && y == 7'd355) || (x == 203 && y == 264) ||
		(x == 7'd67 && y == 7'd637) || (x == 454 && y == 423) || (x == 7'd30 && y == 489) ||
		(x == 7'd321 && y == 7'd346) || (x == 7'd146 && y == 218) || (x == 438 && y == 7'd423) ||
		(x == 7'd263 && y == 7'd281) || (x == 333 && y == 7'd538) || (x == 328 && y == 540) ||
		(x == 56 && y == 7'd273) || (x == 184 && y == 610) || (x == 458 && y == 7'd477) ||
		(x == 7'd574 && y == 7'd557) || (x == 460 && y == 621) || (x == 7'd278 && y == 413) ||
		(x == 7'd41 && y == 7'd261) || (x == 7'd69 && y == 311) || (x == 307 && y == 212) ||
		(x == 7'd210 && y == 7'd567) || (x == 454 && y == 473) || (x == 7'd553 && y == 62) ||
		(x == 7'd396 && y == 7'd625) || (x == 265 && y == 7'd332) || (x == 7'd343 && y == 16) ||
		(x == 7'd455 && y == 535) || (x == 547 && y == 368) || (x == 349 && y == 7'd341) ||
		(x == 7'd251 && y == 7'd312) || (x == 7'd108 && y == 428) || (x == 338 && y == 7'd461) ||
		(x == 7'd486 && y == 7'd366) || (x == 372 && y == 7'd152) || (x == 225 && y == 423) ||
		(x == 381 && y == 571) || (x == 401 && y == 7'd149) || (x == 176 && y == 154) ||
		(x == 573 && y == 7'd240) || (x == 7'd412 && y == 636) || (x == 291 && y == 245) ||
		(x == 7'd422 && y == 621) || (x == 623 && y == 282) || (x == 7'd144 && y == 7'd209) ||
		(x == 7'd228 && y == 332) || (x == 7'd310 && y == 200) || (x == 161 && y == 7'd218) ||
		(x == 604 && y == 413) || (x == 7'd107 && y == 222) || (x == 7'd484 && y == 7'd551) ||
		(x == 611 && y == 583) || (x == 247 && y == 7'd220) || (x == 7'd368 && y == 7'd132) ||
		(x == 7'd388 && y == 7'd561) || (x == 7'd121 && y == 7'd169) || (x == 277 && y == 7'd80) ||
		(x == 7'd250 && y == 7'd597) || (x == 271 && y == 321) || (x == 7'd614 && y == 7'd256) ||
		(x == 7'd599 && y == 7'd619) || (x == 7'd540 && y == 7'd301) || (x == 7'd186 && y == 7'd634) ||
		(x == 7'd445 && y == 7'd66) || (x == 397 && y == 176) || (x == 7'd125 && y == 524) ||
		(x == 7'd220 && y == 7'd142) || (x == 615 && y == 525) || (x == 249 && y == 547) ||
		(x == 7'd542 && y == 7'd84) || (x == 7'd76 && y == 562) || (x == 581 && y == 234) ||
		(x == 386 && y == 310) || (x == 7'd472 && y == 7'd150) || (x == 7'd374 && y == 253) ||
		(x == 7'd631 && y == 7'd56) || (x == 7'd201 && y == 292) || (x == 146 && y == 7'd526) ||
		(x == 287 && y == 548) || (x == 7'd334 && y == 328) || (x == 7'd126 && y == 192) ||
		(x == 560 && y == 7'd106) || (x == 7'd516 && y == 12) || (x == 530 && y == 256) ||
		(x == 7'd23 && y == 204) || (x == 450 && y == 7'd82) || (x == 7'd153 && y == 582) ||
		(x == 476 && y == 7'd168) || (x == 7'd237 && y == 7'd597) || (x == 167 && y == 408) ||
		(x == 7'd249 && y == 7'd611) || (x == 7'd461 && y == 7'd128) || (x == 281 && y == 7'd483) ||
		(x == 7'd240 && y == 7'd251) || (x == 7'd480 && y == 7'd493) || (x == 7'd89 && y == 7'd625) ||
		(x == 7'd284 && y == 105) || (x == 7'd33 && y == 7'd358) || (x == 7'd279 && y == 77) ||
		(x == 347 && y == 169) || (x == 7'd618 && y == 7'd247) || (x == 7'd409 && y == 7'd3) ||
		(x == 7'd474 && y == 7'd375) || (x == 397 && y == 7'd307) || (x == 7'd595 && y == 374) ||
		(x == 7'd452 && y == 7'd133) || (x == 7'd399 && y == 7'd192) || (x == 601 && y == 561) ||
		(x == 7'd499 && y == 476) || (x == 175 && y == 168) || (x == 172 && y == 507) ||
		(x == 7'd337 && y == 7'd513) || (x == 7'd134 && y == 227) || (x == 7'd191 && y == 7'd40) ||
		(x == 402 && y == 7'd367) || (x == 477 && y == 246) || (x == 7'd237 && y == 18) ||
		(x == 7'd186 && y == 7'd402) || (x == 7'd182 && y == 7'd363) || (x == 113 && y == 7'd165) ||
		(x == 632 && y == 185) || (x == 7'd298 && y == 270) || (x == 7'd589 && y == 222) ||
		(x == 7'd547 && y == 316) || (x == 7'd468 && y == 7'd374) || (x == 7'd374 && y == 457) ||
		(x == 415 && y == 512) || (x == 513 && y == 411) || (x == 543 && y == 349) ||
		(x == 153 && y == 312) || (x == 7'd554 && y == 225) || (x == 7'd17 && y == 7'd581) ||
		(x == 7'd262 && y == 7'd198) || (x == 614 && y == 7'd281) || (x == 7'd17 && y == 7'd324) ||
		(x == 7'd419 && y == 7'd469) || (x == 155 && y == 7'd212) || (x == 7'd206 && y == 269) ||
		(x == 366 && y == 315) || (x == 546 && y == 132) || (x == 7'd537 && y == 7'd394) ||
		(x == 445 && y == 7'd271) || (x == 7'd372 && y == 318) || (x == 201 && y == 7'd255) ||
		(x == 7'd485 && y == 539) || (x == 7'd504 && y == 7'd234) || (x == 7'd611 && y == 7'd135) ||
		(x == 7'd435 && y == 577) || (x == 7'd200 && y == 7'd269) || (x == 50 && y == 7'd271) ||
		(x == 7'd42 && y == 640) || (x == 630 && y == 7'd462) || (x == 170 && y == 7'd57) ||
		(x == 245 && y == 7'd246) || (x == 235 && y == 7'd31) || (x == 7'd350 && y == 568) ||
		(x == 625 && y == 509) || (x == 545 && y == 7'd98) || (x == 568 && y == 7'd116) ||
		(x == 279 && y == 441) || (x == 322 && y == 7'd169) || (x == 508 && y == 580) ||
		(x == 558 && y == 7'd390) || (x == 190 && y == 210) || (x == 178 && y == 7'd627) ||
		(x == 7'd297 && y == 7'd341) || (x == 7'd249 && y == 7'd311) || (x == 7'd63 && y == 82) ||
		(x == 544 && y == 7'd69) || (x == 7'd569 && y == 507) || (x == 7'd579 && y == 7'd619) ||
		(x == 379 && y == 431) || (x == 12 && y == 7'd169) || (x == 7'd5 && y == 28) ||
		(x == 134 && y == 7'd368) || (x == 7'd540 && y == 7'd394) || (x == 7'd234 && y == 95) ||
		(x == 7'd363 && y == 7'd626) || (x == 7'd397 && y == 7'd441) || (x == 7'd334 && y == 7'd435) ||
		(x == 295 && y == 7'd159) || (x == 7'd101 && y == 213) || (x == 407 && y == 297) ||
		(x == 7'd615 && y == 7'd104) || (x == 456 && y == 7'd456) || (x == 7'd44 && y == 7'd340) ||
		(x == 7'd99 && y == 295) || (x == 7'd623 && y == 7'd479) || (x == 468 && y == 635) ||
		(x == 514 && y == 7'd47) || (x == 7'd582 && y == 223) || (x == 7'd518 && y == 7'd246) ||
		(x == 7'd59 && y == 7'd223) || (x == 7'd457 && y == 4) || (x == 7'd163 && y == 7'd399) ||
		(x == 231 && y == 7'd165) || (x == 289 && y == 175) || (x == 7'd308 && y == 7'd446) ||
		(x == 130 && y == 637) || (x == 7'd490 && y == 7'd429) || (x == 7'd407 && y == 274) ||
		(x == 7'd123 && y == 7'd409) || (x == 7'd95 && y == 7'd566) || (x == 7'd95 && y == 7'd391) ||
		(x == 340 && y == 148) || (x == 152 && y == 265) || (x == 190 && y == 214) ||
		(x == 7'd96 && y == 389) || (x == 7'd495 && y == 7'd624) || (x == 411 && y == 549) ||
		(x == 7'd225 && y == 7'd363) || (x == 423 && y == 266) || (x == 7'd508 && y == 7'd42) ||
		(x == 7'd426 && y == 468) || (x == 7'd159 && y == 271) || (x == 7'd415 && y == 7'd398) ||
		(x == 543 && y == 373) || (x == 460 && y == 615) || (x == 7'd136 && y == 11) ||
		(x == 7'd323 && y == 470) || (x == 324 && y == 7'd482) || (x == 311 && y == 603) ||
		(x == 597 && y == 454) || (x == 7'd251 && y == 7'd593) || (x == 7'd292 && y == 7'd143) ||
		(x == 7'd274 && y == 274) || (x == 7'd348 && y == 7'd380) || (x == 112 && y == 7'd180) ||
		(x == 597 && y == 362) || (x == 579 && y == 7'd307) || (x == 7'd487 && y == 374) ||
		(x == 565 && y == 7'd604) || (x == 7'd364 && y == 7'd435) || (x == 7'd353 && y == 7'd393) ||
		(x == 7'd280 && y == 501) || (x == 316 && y == 7'd238) || (x == 242 && y == 244) ||
		(x == 7'd191 && y == 7'd619) || (x == 7'd103 && y == 7'd455) || (x == 223 && y == 507) ||
		(x == 7'd200 && y == 7'd566) || (x == 7'd621 && y == 620) || (x == 369 && y == 7'd602) ||
		(x == 231 && y == 475) || (x == 477 && y == 566) || (x == 7'd205 && y == 480) ||
		(x == 7'd434 && y == 464) || (x == 7'd400 && y == 7'd241) || (x == 277 && y == 369) ||
		(x == 7'd217 && y == 7'd496) || (x == 7'd248 && y == 7'd14) || (x == 7'd399 && y == 7'd503) ||
		(x == 7'd387 && y == 7'd488) || (x == 175 && y == 7'd157) || (x == 7'd584 && y == 7'd529) ||
		(x == 390 && y == 403) || (x == 443 && y == 7'd376) || (x == 7'd580 && y == 7'd463) ||
		(x == 7'd610 && y == 7'd549) || (x == 193 && y == 243) || (x == 7'd208 && y == 7'd107) ||
		(x == 221 && y == 7'd132) || (x == 7'd605 && y == 7'd123) || (x == 254 && y == 7'd281) ||
		(x == 7'd576 && y == 212) || (x == 471 && y == 7'd487) || (x == 7'd267 && y == 7'd535) ||
		(x == 272 && y == 282) || (x == 7'd28 && y == 7'd258) || (x == 349 && y == 411) ||
		(x == 7'd275 && y == 7'd410) || (x == 7'd406 && y == 237) || (x == 7'd616 && y == 7'd208) ||
		(x == 7'd364 && y == 7'd515) || (x == 7'd509 && y == 7'd299) || (x == 7'd438 && y == 7'd145) ||
		(x == 259 && y == 493) || (x == 389 && y == 535) || (x == 7'd76 && y == 7'd155) ||
		(x == 7'd516 && y == 7'd560) || (x == 7'd226 && y == 628) || (x == 7'd491 && y == 7'd468) ||
		(x == 318 && y == 7'd528) || (x == 7'd611 && y == 7'd259) || (x == 7'd300 && y == 7'd465) ||
		(x == 7'd181 && y == 519) || (x == 7'd597 && y == 7'd118) || (x == 337 && y == 7'd391) ||
		(x == 579 && y == 136) || (x == 406 && y == 7'd295) || (x == 172 && y == 7'd538) ||
		(x == 7'd160 && y == 7'd399) || (x == 7'd394 && y == 7'd500) || (x == 584 && y == 446) ||
		(x == 550 && y == 399) || (x == 334 && y == 363) || (x == 368 && y == 7'd290) ||
		(x == 7'd95 && y == 477) || (x == 7'd449 && y == 7'd594) || (x == 536 && y == 7'd408) ||
		(x == 7'd92 && y == 419) || (x == 150 && y == 7'd382) || (x == 573 && y == 7'd601) ||
		(x == 514 && y == 7'd441) || (x == 10 && y == 7'd152) || (x == 7'd209 && y == 7'd467) ||
		(x == 7'd608 && y == 7'd361) || (x == 223 && y == 405) || (x == 503 && y == 7'd618) ||
		(x == 7'd97 && y == 258) || (x == 7'd548 && y == 7'd347) || (x == 595 && y == 7'd229) ||
		(x == 7'd220 && y == 564) || (x == 7'd625 && y == 7'd518) || (x == 148 && y == 7'd251) ||
		(x == 7'd616 && y == 7'd132) || (x == 7'd185 && y == 7'd258) || (x == 7'd295 && y == 7'd498) ||
		(x == 7'd388 && y == 242) || (x == 7'd445 && y == 606) || (x == 7'd428 && y == 10) ||
		(x == 7'd85 && y == 107) || (x == 7'd582 && y == 7'd134) || (x == 7'd599 && y == 161) ||
		(x == 7'd207 && y == 28) || (x == 7'd412 && y == 592) || (x == 7'd590 && y == 7'd124) ||
		(x == 301 && y == 7'd609) || (x == 7'd437 && y == 210) || (x == 227 && y == 7'd62) ||
		(x == 364 && y == 7'd479) || (x == 7'd168 && y == 7'd514) || (x == 7'd380 && y == 310) ||
		(x == 7'd443 && y == 100) || (x == 579 && y == 7'd324) || (x == 458 && y == 7'd522) ||
		(x == 7'd626 && y == 7'd577) || (x == 529 && y == 7'd588) || (x == 7'd422 && y == 233) ||
		(x == 269 && y == 7'd467) || (x == 429 && y == 607) || (x == 613 && y == 7'd273) ||
		(x == 7'd292 && y == 253) || (x == 7'd38 && y == 7'd489) || (x == 292 && y == 421) ||
		(x == 7'd577 && y == 7'd572) || (x == 7'd526 && y == 146) || (x == 7'd94 && y == 282) ||
		(x == 7'd189 && y == 7'd85) || (x == 7'd229 && y == 7'd484) || (x == 7'd220 && y == 376) ||
		(x == 160 && y == 7'd128) || (x == 7'd70 && y == 7'd566) || (x == 7'd582 && y == 7'd110) ||
		(x == 7'd58 && y == 7'd512) || (x == 7'd347 && y == 7'd527) || (x == 42 && y == 7'd397) ||
		(x == 124 && y == 7'd300) || (x == 7'd639 && y == 7'd341) || (x == 272 && y == 7'd613) ||
		(x == 60 && y == 7'd247) || (x == 7'd191 && y == 7'd450) || (x == 7'd603 && y == 7'd395) ||
		(x == 7'd377 && y == 7'd510) || (x == 7'd543 && y == 7'd508) || (x == 7'd482 && y == 39) ||
		(x == 7'd520 && y == 7'd419) || (x == 7'd296 && y == 7'd131) || (x == 7'd537 && y == 339) ||
		(x == 7'd594 && y == 7'd601) || (x == 93 && y == 7'd124) || (x == 537 && y == 381) ||
		(x == 7'd309 && y == 7'd619) || (x == 7'd311 && y == 7'd613) || (x == 521 && y == 185) ||
		(x == 7'd590 && y == 594) || (x == 7'd419 && y == 7'd0) || (x == 7'd204 && y == 7'd426) ||
		(x == 7'd189 && y == 7'd373) || (x == 7'd618 && y == 7'd243) || (x == 7'd164 && y == 582) ||
		(x == 515 && y == 7'd608) || (x == 7'd150 && y == 393) || (x == 7'd395 && y == 274) ||
		(x == 7'd257 && y == 376) || (x == 7'd595 && y == 7'd368) || (x == 7'd371 && y == 7'd585) ||
		(x == 7'd74 && y == 314) || (x == 7'd597 && y == 7'd601) || (x == 613 && y == 135) ||
		(x == 479 && y == 7'd413) || (x == 7'd539 && y == 371) || (x == 7'd265 && y == 7'd477) ||
		(x == 498 && y == 129) || (x == 7'd123 && y == 7'd121) || (x == 7'd388 && y == 5) ||
		(x == 521 && y == 7'd25) || (x == 174 && y == 7'd579) || (x == 618 && y == 7'd460) ||
		(x == 18 && y == 7'd268) || (x == 7'd437 && y == 531) || (x == 7'd625 && y == 7'd271) ||
		(x == 7'd320 && y == 626) || (x == 39 && y == 7'd238) || (x == 7'd507 && y == 441) ||
		(x == 7'd203 && y == 7'd259) || (x == 549 && y == 7'd48) || (x == 263 && y == 297) ||
		(x == 7'd171 && y == 345) || (x == 7'd626 && y == 7'd271) || (x == 7'd398 && y == 7'd532) ||
		(x == 7'd619 && y == 22) || (x == 7'd190 && y == 7'd91) || (x == 28 && y == 7'd161) ||
		(x == 7'd2 && y == 459) || (x == 181 && y == 287) || (x == 190 && y == 7'd420) ||
		(x == 441 && y == 7'd241) || (x == 7'd50 && y == 420) || (x == 578 && y == 223) ||
		(x == 7'd589 && y == 7'd50) || (x == 7'd340 && y == 7'd340) || (x == 396 && y == 7'd640) ||
		(x == 7'd210 && y == 7'd114) || (x == 7'd226 && y == 7'd388) || (x == 460 && y == 507) ||
		(x == 7'd271 && y == 7'd529) || (x == 589 && y == 7'd223) || (x == 480 && y == 507) ||
		(x == 7'd123 && y == 209) || (x == 7'd609 && y == 7'd8) || (x == 403 && y == 7'd103) ||
		(x == 7'd549 && y == 7'd294) || (x == 7'd146 && y == 7'd415) || (x == 388 && y == 7'd241) ||
		(x == 198 && y == 253) || (x == 7'd434 && y == 16) || (x == 178 && y == 7'd617) ||
		(x == 7'd285 && y == 7'd398) || (x == 7'd573 && y == 252) || (x == 7'd435 && y == 7'd386) ||
		(x == 324 && y == 7'd317) || (x == 484 && y == 7'd626) || (x == 7'd350 && y == 7'd369) ||
		(x == 578 && y == 341) || (x == 7'd599 && y == 234) || (x == 7'd372 && y == 7'd477) ||
		(x == 7'd499 && y == 7'd546) || (x == 7'd253 && y == 7'd424) || (x == 7'd556 && y == 7'd637) ||
		(x == 19 && y == 7'd173) || (x == 7'd73 && y == 199) || (x == 7'd358 && y == 7'd458) ||
		(x == 7'd303 && y == 156) || (x == 7'd214 && y == 7'd245) || (x == 7'd132 && y == 7'd47) ||
		(x == 271 && y == 7'd538) || (x == 7'd530 && y == 7'd555) || (x == 345 && y == 7'd207) ||
		(x == 229 && y == 498) || (x == 515 && y == 591) || (x == 616 && y == 7'd82) ||
		(x == 7'd131 && y == 7'd391) || (x == 339 && y == 338) || (x == 7'd634 && y == 610) ||
		(x == 7'd328 && y == 357) || (x == 186 && y == 163) || (x == 365 && y == 7'd134) ||
		(x == 7'd616 && y == 587) || (x == 7'd64 && y == 7'd264) || (x == 7'd328 && y == 7'd508) ||
		(x == 7'd369 && y == 7'd500) || (x == 451 && y == 7'd282) || (x == 10 && y == 7'd269) ||
		(x == 7'd367 && y == 7'd271) || (x == 157 && y == 429) || (x == 292 && y == 351) ||
		(x == 547 && y == 359) || (x == 7'd358 && y == 7'd507) || (x == 7'd368 && y == 7'd453) ||
		(x == 534 && y == 7'd178) || (x == 7'd137 && y == 7'd497) || (x == 7'd312 && y == 7'd209) ||
		(x == 284 && y == 285) || (x == 7'd206 && y == 629) || (x == 7'd620 && y == 7'd431) ||
		(x == 7'd536 && y == 7'd363) || (x == 370 && y == 463) || (x == 538 && y == 195) ||
		(x == 362 && y == 304) || (x == 526 && y == 7'd83) || (x == 7'd387 && y == 7'd612) ||
		(x == 7'd579 && y == 133) || (x == 7'd239 && y == 7'd130) || (x == 7'd368 && y == 7'd506) ||
		(x == 209 && y == 207) || (x == 7'd559 && y == 622) || (x == 220 && y == 7'd60) ||
		(x == 7'd283 && y == 7'd522) || (x == 7'd421 && y == 7'd37) || (x == 7'd439 && y == 277) ||
		(x == 7'd183 && y == 227) || (x == 7'd136 && y == 7'd288) || (x == 7'd398 && y == 38) ||
		(x == 580 && y == 148) || (x == 276 && y == 190) || (x == 582 && y == 7'd529) ||
		(x == 7'd413 && y == 7'd586) || (x == 7'd443 && y == 7'd491) || (x == 541 && y == 356) ||
		(x == 329 && y == 489) || (x == 7'd494 && y == 7'd518) || (x == 7'd15 && y == 7'd186) ||
		(x == 7'd59 && y == 7'd342) || (x == 258 && y == 320) || (x == 7'd472 && y == 7'd216) ||
		(x == 7'd183 && y == 7'd460) || (x == 7'd182 && y == 7'd496) || (x == 34 && y == 7'd502) ||
		(x == 640 && y == 444) || (x == 7'd459 && y == 7'd179) || (x == 491 && y == 376) ||
		(x == 7'd170 && y == 245) || (x == 7'd89 && y == 590) || (x == 7'd350 && y == 608) ||
		(x == 7'd433 && y == 7'd389) || (x == 161 && y == 7'd253) || (x == 7'd35 && y == 7'd473) ||
		(x == 7'd269 && y == 7'd83) || (x == 132 && y == 353) || (x == 251 && y == 231) ||
		(x == 135 && y == 7'd101) || (x == 7'd60 && y == 7'd633) || (x == 7'd391 && y == 117) ||
		(x == 248 && y == 7'd414) || (x == 220 && y == 7'd530) || (x == 132 && y == 7'd153) ||
		(x == 7'd530 && y == 82) || (x == 7'd637 && y == 7'd565) || (x == 421 && y == 7'd620) ||
		(x == 123 && y == 7'd424) || (x == 7'd460 && y == 196) || (x == 7'd370 && y == 7'd494) ||
		(x == 7'd342 && y == 489) || (x == 7'd228 && y == 183) || (x == 32 && y == 117) ||
		(x == 214 && y == 412) || (x == 7'd106 && y == 117) || (x == 438 && y == 7'd513) ||
		(x == 7'd286 && y == 380) || (x == 379 && y == 429) || (x == 7'd189 && y == 7'd344) ||
		(x == 7'd397 && y == 191) || (x == 473 && y == 7'd404) || (x == 219 && y == 507) ||
		(x == 522 && y == 598) || (x == 7'd365 && y == 7'd24) || (x == 7'd517 && y == 7'd434) ||
		(x == 318 && y == 411) || (x == 8 && y == 7'd68) || (x == 391 && y == 7'd136) ||
		(x == 7'd390 && y == 7'd631) || (x == 7'd624 && y == 7'd504) || (x == 7'd578 && y == 63) ||
		(x == 7'd262 && y == 7'd618) || (x == 279 && y == 465) || (x == 7'd602 && y == 140) ||
		(x == 7'd108 && y == 7'd610) || (x == 7'd34 && y == 565) || (x == 527 && y == 7'd561) ||
		(x == 7'd631 && y == 600) || (x == 160 && y == 344) || (x == 159 && y == 7'd178) ||
		(x == 7'd613 && y == 343) || (x == 7'd183 && y == 483) || (x == 7'd445 && y == 7'd158) ||
		(x == 7'd117 && y == 7'd330) || (x == 7'd358 && y == 7'd411) || (x == 115 && y == 7'd454) ||
		(x == 52 && y == 7'd532) || (x == 505 && y == 7'd198) || (x == 7'd143 && y == 7'd367) ||
		(x == 7'd230 && y == 221) || (x == 7'd310 && y == 7'd274) || (x == 7'd575 && y == 7'd264) ||
		(x == 7'd521 && y == 581) || (x == 155 && y == 7'd472) || (x == 7'd128 && y == 454) ||
		(x == 7'd527 && y == 7'd191) || (x == 7'd15 && y == 184) || (x == 486 && y == 7'd235) ||
		(x == 587 && y == 7'd359) || (x == 632 && y == 373) || (x == 7'd208 && y == 7'd75) ||
		(x == 161 && y == 7'd341) || (x == 7'd421 && y == 132) || (x == 7'd534 && y == 7'd122) ||
		(x == 115 && y == 7'd584) || (x == 7'd69 && y == 354) || (x == 334 && y == 142) ||
		(x == 564 && y == 7'd282) || (x == 7'd267 && y == 7'd334) || (x == 7'd289 && y == 7'd68) ||
		(x == 7'd275 && y == 7'd515) || (x == 11 && y == 7'd291) || (x == 371 && y == 7'd124) ||
		(x == 412 && y == 7'd28) || (x == 7'd311 && y == 7'd402) || (x == 7'd551 && y == 340) ||
		(x == 7'd396 && y == 279) || (x == 7'd381 && y == 243) || (x == 7'd35 && y == 580) ||
		(x == 7'd471 && y == 3) || (x == 51 && y == 7'd512) || (x == 7'd337 && y == 7'd87) ||
		(x == 7'd157 && y == 433) || (x == 7'd634 && y == 7'd530) || (x == 204 && y == 166) ||
		(x == 205 && y == 134) || (x == 7'd150 && y == 575) || (x == 110 && y == 7'd378) ||
		(x == 392 && y == 7'd32) || (x == 7'd579 && y == 7'd175) || (x == 546 && y == 133) ||
		(x == 464 && y == 495) || (x == 7'd458 && y == 7'd617) || (x == 486 && y == 178) ||
		(x == 561 && y == 162) || (x == 187 && y == 245) || (x == 7'd336 && y == 7'd336) ||
		(x == 7'd346 && y == 85) || (x == 560 && y == 455) || (x == 7'd52 && y == 294) ||
		(x == 7'd193 && y == 7'd201) || (x == 7'd347 && y == 152) || (x == 7'd225 && y == 7'd15) ||
		(x == 381 && y == 240) || (x == 7'd13 && y == 7'd499) || (x == 7'd527 && y == 7'd440) ||
		(x == 7'd27 && y == 36) || (x == 154 && y == 544) || (x == 7'd264 && y == 7'd187) ||
		(x == 316 && y == 193) || (x == 476 && y == 7'd359) || (x == 7'd8 && y == 92) ||
		(x == 7'd577 && y == 235) || (x == 552 && y == 599) || (x == 7'd524 && y == 572) ||
		(x == 311 && y == 7'd77) || (x == 7'd217 && y == 7'd503) || (x == 7'd342 && y == 323) ||
		(x == 422 && y == 7'd196) || (x == 7'd150 && y == 7'd583) || (x == 187 && y == 156) ||
		(x == 7'd595 && y == 7'd313) || (x == 7'd431 && y == 171) || (x == 507 && y == 7'd244) ||
		(x == 229 && y == 7'd350) || (x == 7'd539 && y == 7'd308) || (x == 7'd260 && y == 102) ||
		(x == 7'd219 && y == 7'd401) || (x == 300 && y == 537) || (x == 7'd371 && y == 160) ||
		(x == 7'd331 && y == 7'd147) || (x == 7'd238 && y == 7'd300) || (x == 7'd505 && y == 7'd586) ||
		(x == 619 && y == 7'd423) || (x == 556 && y == 7'd158) || (x == 7'd331 && y == 7'd553) ||
		(x == 423 && y == 7'd619) || (x == 411 && y == 474) || (x == 7'd589 && y == 7'd381) ||
		(x == 7'd56 && y == 207) || (x == 7'd451 && y == 7'd497) || (x == 7'd464 && y == 281) ||
		(x == 7'd154 && y == 7'd265) || (x == 468 && y == 7'd511) || (x == 7'd616 && y == 76) ||
		(x == 7'd430 && y == 410) || (x == 7'd261 && y == 7'd477) || (x == 7'd242 && y == 298) ||
		(x == 7'd294 && y == 7'd457) || (x == 7'd192 && y == 371) || (x == 7'd377 && y == 7'd204) ||
		(x == 154 && y == 303) || (x == 477 && y == 7'd125) || (x == 7'd571 && y == 7'd2) ||
		(x == 581 && y == 277) || (x == 581 && y == 7'd637) || (x == 238 && y == 526) ||
		(x == 7'd564 && y == 7'd433) || (x == 7'd100 && y == 602) || (x == 7'd617 && y == 261) ||
		(x == 355 && y == 7'd520) || (x == 7'd546 && y == 7'd578) || (x == 7'd560 && y == 7'd208) ||
		(x == 321 && y == 157) || (x == 184 && y == 7'd492) || (x == 7'd186 && y == 7'd613) ||
		(x == 7'd155 && y == 328) || (x == 7'd570 && y == 577) || (x == 256 && y == 412) ||
		(x == 627 && y == 7'd270) || (x == 7'd291 && y == 7'd64) || (x == 7'd441 && y == 7'd147) ||
		(x == 256 && y == 7'd89) || (x == 405 && y == 371) || (x == 7'd157 && y == 441) ||
		(x == 7'd632 && y == 7'd191) || (x == 7'd453 && y == 7'd617) || (x == 7'd329 && y == 7'd552) ||
		(x == 7'd374 && y == 505) || (x == 7'd509 && y == 7'd306) || (x == 437 && y == 7'd265) ||
		(x == 7'd564 && y == 7'd76) || (x == 7'd147 && y == 7'd308) || (x == 58 && y == 7'd455) ||
		(x == 7'd381 && y == 7'd629) || (x == 93 && y == 7'd293) || (x == 357 && y == 7'd369) ||
		(x == 88 && y == 7'd157) || (x == 572 && y == 549) || (x == 7'd273 && y == 7'd469) ||
		(x == 7'd603 && y == 8) || (x == 7'd61 && y == 7'd554) || (x == 575 && y == 7'd525) ||
		(x == 7'd508 && y == 7'd307) || (x == 7'd234 && y == 7'd472) || (x == 163 && y == 7'd622) ||
		(x == 545 && y == 7'd486) || (x == 7'd374 && y == 7'd589) || (x == 396 && y == 600) ||
		(x == 390 && y == 7'd46) || (x == 7'd349 && y == 402) || (x == 7'd85 && y == 250) ||
		(x == 7'd229 && y == 7'd260) || (x == 7'd200 && y == 7'd412) || (x == 261 && y == 154) ||
		(x == 260 && y == 7'd628) || (x == 281 && y == 7'd211) || (x == 555 && y == 136) ||
		(x == 7'd306 && y == 377) || (x == 306 && y == 7'd457) || (x == 135 && y == 7'd394) ||
		(x == 7'd394 && y == 7'd22) || (x == 257 && y == 576) || (x == 202 && y == 7'd362) ||
		(x == 7'd291 && y == 7'd528) || (x == 7'd66 && y == 335) || (x == 19 && y == 33) ||
		(x == 7'd250 && y == 7'd299) || (x == 7'd164 && y == 606) || (x == 7'd603 && y == 169) ||
		(x == 7'd517 && y == 7'd362) || (x == 7'd521 && y == 7'd185) || (x == 565 && y == 7'd449) ||
		(x == 7'd68 && y == 73) || (x == 499 && y == 7'd383) || (x == 7'd142 && y == 598) ||
		(x == 7'd377 && y == 16) || (x == 525 && y == 7'd61) || (x == 7'd380 && y == 476) ||
		(x == 7'd309 && y == 7'd513) || (x == 352 && y == 260) || (x == 580 && y == 7'd407) ||
		(x == 7'd187 && y == 141) || (x == 7'd160 && y == 7'd196) || (x == 7'd420 && y == 7'd114) ||
		(x == 539 && y == 7'd347) || (x == 119 && y == 7'd611) || (x == 7'd144 && y == 7'd500) ||
		(x == 321 && y == 164) || (x == 615 && y == 7'd22) || (x == 199 && y == 7'd412) ||
		(x == 7'd37 && y == 367) || (x == 7'd68 && y == 241) || (x == 440 && y == 141) ||
		(x == 7'd199 && y == 7'd185) || (x == 7'd423 && y == 176) || (x == 7'd525 && y == 182) ||
		(x == 7'd40 && y == 411) || (x == 7'd524 && y == 81) || (x == 7'd391 && y == 168) ||
		(x == 212 && y == 7'd342) || (x == 402 && y == 508) || (x == 7'd253 && y == 203) ||
		(x == 7'd92 && y == 7'd50) || (x == 7'd210 && y == 7'd468) || (x == 349 && y == 470) ||
		(x == 7'd123 && y == 7'd19) || (x == 151 && y == 419) || (x == 7'd373 && y == 7'd624) ||
		(x == 378 && y == 561) || (x == 7'd404 && y == 429) || (x == 4 && y == 7'd567) ||
		(x == 246 && y == 7'd113) || (x == 7'd341 && y == 7'd592) || (x == 7'd449 && y == 7'd192) ||
		(x == 7'd635 && y == 7'd569) || (x == 7'd607 && y == 221) || (x == 7'd493 && y == 7'd532) ||
		(x == 114 && y == 7'd71) || (x == 7'd443 && y == 7'd324) || (x == 281 && y == 331) ||
		(x == 254 && y == 7'd184) || (x == 393 && y == 7'd192) || (x == 10 && y == 7'd514) ||
		(x == 636 && y == 7'd328) || (x == 7'd404 && y == 7'd173) || (x == 574 && y == 7'd387) ||
		(x == 7'd449 && y == 7'd595) || (x == 7'd391 && y == 7'd524) || (x == 7'd414 && y == 7'd17) ||
		(x == 420 && y == 220) || (x == 129 && y == 7'd122) || (x == 554 && y == 7'd275) ||
		(x == 7'd392 && y == 7'd623) || (x == 7'd392 && y == 7'd276) || (x == 7'd53 && y == 611) ||
		(x == 7'd372 && y == 7'd287) || (x == 13 && y == 7'd602) || (x == 640 && y == 7'd601) ||
		(x == 7'd276 && y == 596) || (x == 594 && y == 567) || (x == 7'd355 && y == 394) ||
		(x == 496 && y == 7'd495) || (x == 7'd198 && y == 7'd258) || (x == 263 && y == 552) ||
		(x == 7'd428 && y == 7'd95) || (x == 305 && y == 7'd419) || (x == 512 && y == 7'd532) ||
		(x == 7'd117 && y == 620) || (x == 9 && y == 7'd296) || (x == 7'd123 && y == 144) ||
		(x == 7'd133 && y == 7'd525) || (x == 7'd161 && y == 557) || (x == 162 && y == 512) ||
		(x == 7'd595 && y == 7'd445) || (x == 7'd346 && y == 7'd529) || (x == 7'd391 && y == 300) ||
		(x == 366 && y == 7'd496) || (x == 7'd460 && y == 575) || (x == 503 && y == 481) ||
		(x == 7'd384 && y == 192) || (x == 7'd606 && y == 107) || (x == 7'd200 && y == 7'd331) ||
		(x == 145 && y == 390) || (x == 528 && y == 7'd61) || (x == 257 && y == 234) ||
		(x == 7'd612 && y == 7'd258) || (x == 196 && y == 496) || (x == 165 && y == 7'd591) ||
		(x == 587 && y == 7'd588) || (x == 322 && y == 144) || (x == 7'd425 && y == 7'd170) ||
		(x == 7'd368 && y == 217) || (x == 407 && y == 243) || (x == 591 && y == 536) ||
		(x == 620 && y == 145) || (x == 7'd45 && y == 7'd265) || (x == 7'd496 && y == 7'd439) ||
		(x == 477 && y == 624) || (x == 7'd387 && y == 7'd479) || (x == 215 && y == 7'd550) ||
		(x == 307 && y == 586) || (x == 617 && y == 7'd4) || (x == 7'd574 && y == 430) ||
		(x == 7'd133 && y == 7'd508) || (x == 326 && y == 321) || (x == 7'd230 && y == 7'd81) ||
		(x == 7'd131 && y == 97) || (x == 230 && y == 616) || (x == 503 && y == 281) ||
		(x == 163 && y == 248) || (x == 7'd629 && y == 7'd602) || (x == 533 && y == 7'd176) ||
		(x == 395 && y == 7'd111) || (x == 7'd263 && y == 501) || (x == 7'd129 && y == 529) ||
		(x == 7'd284 && y == 7'd253) || (x == 148 && y == 471) || (x == 7'd623 && y == 7'd513) ||
		(x == 7'd39 && y == 486) || (x == 585 && y == 287) || (x == 200 && y == 317) ||
		(x == 7'd562 && y == 285) || (x == 179 && y == 214) || (x == 7'd48 && y == 497) ||
		(x == 7'd483 && y == 412) || (x == 444 && y == 7'd165) || (x == 7'd575 && y == 65) ||
		(x == 7'd203 && y == 7'd180) || (x == 7'd249 && y == 7'd509) || (x == 452 && y == 172) ||
		(x == 139 && y == 7'd360) || (x == 216 && y == 326) || (x == 214 && y == 7'd630) ||
		(x == 393 && y == 343) || (x == 7'd273 && y == 7'd528) || (x == 7'd469 && y == 7'd52) ||
		(x == 7'd526 && y == 7'd320) || (x == 7'd379 && y == 7'd132) || (x == 7'd586 && y == 357) ||
		(x == 188 && y == 407) || (x == 130 && y == 526) || (x == 7'd337 && y == 7'd356) ||
		(x == 7'd357 && y == 7'd591) || (x == 336 && y == 7'd104) || (x == 7'd195 && y == 7'd302) ||
		(x == 7'd251 && y == 220) || (x == 7'd7 && y == 7'd278) || (x == 127 && y == 7'd204) ||
		(x == 7'd366 && y == 426) || (x == 504 && y == 7'd20) || (x == 7'd284 && y == 7'd140) ||
		(x == 7'd441 && y == 346) || (x == 603 && y == 7'd362) || (x == 7'd197 && y == 7'd358) ||
		(x == 7'd573 && y == 7'd105) || (x == 227 && y == 208) || (x == 397 && y == 7'd412) ||
		(x == 283 && y == 7'd408) || (x == 7'd586 && y == 146) || (x == 7'd512 && y == 278) ||
		(x == 42 && y == 7'd263) || (x == 14 && y == 7'd419) || (x == 7'd631 && y == 7'd36) ||
		(x == 7'd40 && y == 205) || (x == 7'd82 && y == 7'd376) || (x == 283 && y == 7'd637) ||
		(x == 7'd255 && y == 485) || (x == 7'd365 && y == 53) || (x == 569 && y == 7'd83) ||
		(x == 7'd581 && y == 322) || (x == 135 && y == 259) || (x == 495 && y == 376) ||
		(x == 7'd394 && y == 7'd368) || (x == 7'd485 && y == 562) || (x == 355 && y == 7'd614) ||
		(x == 639 && y == 7'd527) || (x == 40 && y == 7'd339) || (x == 7'd496 && y == 7'd285) ||
		(x == 7'd414 && y == 410) || (x == 7'd436 && y == 7'd529) || (x == 455 && y == 200) ||
		(x == 7'd499 && y == 272) || (x == 7'd66 && y == 7'd424) || (x == 449 && y == 486) ||
		(x == 7'd375 && y == 37) || (x == 529 && y == 7'd528) || (x == 7'd214 && y == 7'd273) ||
		(x == 7'd358 && y == 105) || (x == 7'd386 && y == 7'd615) || (x == 402 && y == 578) ||
		(x == 383 && y == 7'd139) || (x == 7'd502 && y == 535) || (x == 7'd380 && y == 274) ||
		(x == 7'd357 && y == 7'd517) || (x == 7'd572 && y == 260) || (x == 7'd601 && y == 528) ||
		(x == 211 && y == 208) || (x == 7'd267 && y == 440) || (x == 7'd549 && y == 7'd260) ||
		(x == 7'd593 && y == 7'd355) || (x == 7'd408 && y == 466) || (x == 7'd436 && y == 7'd612) ||
		(x == 7'd456 && y == 112) || (x == 7'd519 && y == 602) || (x == 264 && y == 7'd170) ||
		(x == 7'd473 && y == 477) || (x == 7'd600 && y == 7'd626) || (x == 7'd210 && y == 7'd501) ||
		(x == 241 && y == 461) || (x == 476 && y == 401) || (x == 7'd596 && y == 182) ||
		(x == 161 && y == 7'd550) || (x == 7'd398 && y == 519) || (x == 396 && y == 339) ||
		(x == 7'd386 && y == 7'd481) || (x == 7'd142 && y == 364) || (x == 197 && y == 534) ||
		(x == 500 && y == 7'd489) || (x == 7'd508 && y == 104) || (x == 7'd166 && y == 7'd246) ||
		(x == 7'd247 && y == 7'd100) || (x == 7'd560 && y == 179) || (x == 151 && y == 254) ||
		(x == 7'd414 && y == 7'd578) || (x == 259 && y == 7'd593) || (x == 7'd473 && y == 7'd378) ||
		(x == 7'd137 && y == 7'd336) || (x == 382 && y == 249) || (x == 518 && y == 7'd280) ||
		(x == 371 && y == 7'd202) || (x == 7'd590 && y == 7'd275) || (x == 7'd570 && y == 7'd507) ||
		(x == 7'd156 && y == 7'd585) || (x == 176 && y == 237) || (x == 222 && y == 518) ||
		(x == 7'd447 && y == 7'd576) || (x == 7'd494 && y == 627) || (x == 7'd472 && y == 7'd271) ||
		(x == 581 && y == 7'd595) || (x == 7'd58 && y == 618) || (x == 7'd531 && y == 7'd128) ||
		(x == 7'd245 && y == 7'd70) || (x == 7'd547 && y == 7'd83) || (x == 187 && y == 431) ||
		(x == 7'd458 && y == 347) || (x == 204 && y == 460) || (x == 436 && y == 7'd603) ||
		(x == 7'd258 && y == 7'd382) || (x == 7'd211 && y == 119) || (x == 351 && y == 361) ||
		(x == 483 && y == 176) || (x == 7'd95 && y == 375) || (x == 7'd631 && y == 7'd595) ||
		(x == 173 && y == 7'd299) || (x == 7'd133 && y == 198) || (x == 336 && y == 7'd370) ||
		(x == 7'd11 && y == 450) || (x == 7'd587 && y == 395) || (x == 7'd1 && y == 471) ||
		(x == 371 && y == 7'd26) || (x == 287 && y == 7'd25) || (x == 7'd591 && y == 263) ||
		(x == 365 && y == 245) || (x == 7'd415 && y == 7'd375) || (x == 7'd53 && y == 244) ||
		(x == 7'd142 && y == 7'd145) || (x == 6 && y == 7'd534) || (x == 7'd337 && y == 7'd240) ||
		(x == 401 && y == 7'd625) || (x == 496 && y == 7'd410) || (x == 7'd338 && y == 7'd512) ||
		(x == 7'd522 && y == 7'd550) || (x == 7'd290 && y == 7'd212) || (x == 433 && y == 533) ||
		(x == 476 && y == 7'd378) || (x == 596 && y == 537) || (x == 562 && y == 7'd293) ||
		(x == 591 && y == 509) || (x == 7'd521 && y == 7'd142) || (x == 496 && y == 7'd409) ||
		(x == 7'd218 && y == 7'd634) || (x == 7'd467 && y == 197) || (x == 7'd497 && y == 350) ||
		(x == 620 && y == 7'd187) || (x == 178 && y == 142) || (x == 7'd370 && y == 7'd242) ||
		(x == 607 && y == 157) || (x == 7'd130 && y == 7'd395) || (x == 273 && y == 7'd437) ||
		(x == 106 && y == 7'd242) || (x == 232 && y == 322) || (x == 292 && y == 429) ||
		(x == 169 && y == 309) || (x == 7'd98 && y == 7'd183) || (x == 383 && y == 247) ||
		(x == 7'd267 && y == 7'd514) || (x == 7'd329 && y == 7'd105) || (x == 7'd504 && y == 7'd225) ||
		(x == 570 && y == 7'd493) || (x == 7'd22 && y == 355) || (x == 7'd311 && y == 7'd327) ||
		(x == 7'd131 && y == 103) || (x == 7'd370 && y == 7'd221) || (x == 639 && y == 7'd142) ||
		(x == 7'd604 && y == 7'd263) || (x == 34 && y == 7'd629) || (x == 7'd258 && y == 7'd224) ||
		(x == 227 && y == 599) || (x == 7'd567 && y == 582) || (x == 7'd156 && y == 7'd174) ||
		(x == 7'd56 && y == 586) || (x == 350 && y == 7'd251) || (x == 252 && y == 7'd393) ||
		(x == 7'd275 && y == 7'd441) || (x == 7'd120 && y == 7'd287) || (x == 7'd476 && y == 502) ||
		(x == 7'd610 && y == 7) || (x == 591 && y == 326) || (x == 6 && y == 7'd636) ||
		(x == 72 && y == 7'd307) || (x == 7'd568 && y == 7'd467) || (x == 7'd144 && y == 7'd579) ||
		(x == 7'd517 && y == 7'd324) || (x == 271 && y == 7'd134) || (x == 219 && y == 7'd387) ||
		(x == 493 && y == 7'd320) || (x == 582 && y == 7'd339) || (x == 139 && y == 294) ||
		(x == 318 && y == 345) || (x == 7'd520 && y == 7'd401) || (x == 601 && y == 371) ||
		(x == 61 && y == 4) || (x == 7'd381 && y == 7'd529) || (x == 7'd408 && y == 7'd635) ||
		(x == 449 && y == 7'd10) || (x == 239 && y == 388) || (x == 7'd534 && y == 7'd521) ||
		(x == 425 && y == 7'd626) || (x == 300 && y == 540) || (x == 7'd424 && y == 7'd37) ||
		(x == 7'd220 && y == 7'd396) || (x == 11 && y == 7'd90) || (x == 7'd606 && y == 7'd199) ||
		(x == 7'd92 && y == 489) || (x == 7'd391 && y == 313) || (x == 585 && y == 7'd303) ||
		(x == 7'd422 && y == 248) || (x == 406 && y == 7'd189) || (x == 7'd562 && y == 7'd446) ||
		(x == 7'd48 && y == 7'd517) || (x == 455 && y == 184) || (x == 187 && y == 150) ||
		(x == 7'd603 && y == 7'd548) || (x == 431 && y == 7'd96) || (x == 244 && y == 302) ||
		(x == 7'd368 && y == 547) || (x == 7'd160 && y == 7'd619) || (x == 566 && y == 190) ||
		(x == 7'd194 && y == 7'd268) || (x == 7'd150 && y == 120) || (x == 7'd595 && y == 385) ||
		(x == 7'd617 && y == 7'd376) || (x == 628 && y == 315) || (x == 7'd425 && y == 387) ||
		(x == 140 && y == 7'd10) || (x == 7'd218 && y == 429) || (x == 499 && y == 622) ||
		(x == 286 && y == 219) || (x == 7'd280 && y == 327) || (x == 7'd184 && y == 315) ||
		(x == 7'd355 && y == 252) || (x == 7'd464 && y == 7'd489) || (x == 149 && y == 7'd165) ||
		(x == 121 && y == 7'd136) || (x == 7'd421 && y == 475) || (x == 405 && y == 7'd554) ||
		(x == 7'd233 && y == 357) || (x == 129 && y == 7'd314) || (x == 7'd520 && y == 7'd335) ||
		(x == 7'd334 && y == 7'd333) || (x == 261 && y == 7'd70) || (x == 7'd563 && y == 7'd274) ||
		(x == 526 && y == 598) || (x == 187 && y == 552) || (x == 7'd614 && y == 7'd180) ||
		(x == 7'd492 && y == 26) || (x == 608 && y == 599) || (x == 7'd91 && y == 7'd494) ||
		(x == 7'd349 && y == 7'd638) || (x == 467 && y == 7'd561) || (x == 511 && y == 477) ||
		(x == 7'd217 && y == 7'd305) || (x == 220 && y == 365) || (x == 7'd243 && y == 97) ||
		(x == 9 && y == 7'd568) || (x == 7'd250 && y == 7'd635) || (x == 7'd175 && y == 7'd134) ||
		(x == 367 && y == 400) || (x == 7'd420 && y == 7'd387) || (x == 7'd46 && y == 414) ||
		(x == 195 && y == 461) || (x == 140 && y == 7'd230) || (x == 558 && y == 7'd314) ||
		(x == 7'd374 && y == 402) || (x == 7'd23 && y == 7'd207) || (x == 7'd246 && y == 7'd395) ||
		(x == 7'd484 && y == 383) || (x == 7'd357 && y == 424) || (x == 346 && y == 7'd519) ||
		(x == 7'd80 && y == 399) || (x == 224 && y == 574) || (x == 7'd155 && y == 7'd524) ||
		(x == 472 && y == 414) || (x == 7'd278 && y == 7'd560) || (x == 7'd29 && y == 7'd94) ||
		(x == 180 && y == 594) || (x == 7'd466 && y == 7'd62) || (x == 216 && y == 171) ||
		(x == 7'd24 && y == 7'd435) || (x == 7'd118 && y == 7'd295) || (x == 637 && y == 7'd219) ||
		(x == 142 && y == 489) || (x == 7'd409 && y == 7'd132) || (x == 7'd400 && y == 601) ||
		(x == 194 && y == 293) || (x == 7'd48 && y == 371) || (x == 8 && y == 7'd496) ||
		(x == 7'd39 && y == 7'd375) || (x == 7'd144 && y == 7'd297) || (x == 419 && y == 7'd116) ||
		(x == 7'd374 && y == 7'd252) || (x == 7'd155 && y == 7'd226) || (x == 7'd527 && y == 573) ||
		(x == 466 && y == 590) || (x == 278 && y == 380) || (x == 5 && y == 7'd620) ||
		(x == 7'd253 && y == 7'd389) || (x == 7'd52 && y == 546) || (x == 7'd174 && y == 7'd393) ||
		(x == 7'd264 && y == 7'd389) || (x == 196 && y == 7'd510) || (x == 7'd327 && y == 7'd254) ||
		(x == 7'd372 && y == 7'd188) || (x == 558 && y == 373) || (x == 7'd331 && y == 189) ||
		(x == 7'd105 && y == 7'd77) || (x == 123 && y == 7'd555) || (x == 7'd293 && y == 561) ||
		(x == 7'd28 && y == 151) || (x == 632 && y == 7'd520) || (x == 514 && y == 268) ||
		(x == 7'd55 && y == 7'd593) || (x == 295 && y == 7'd278) || (x == 7'd87 && y == 7'd158) ||
		(x == 150 && y == 7'd502) || (x == 7'd35 && y == 7'd130) || (x == 474 && y == 7'd144) ||
		(x == 7'd247 && y == 7'd251) || (x == 306 && y == 7'd510) || (x == 7'd215 && y == 424) ||
		(x == 7'd403 && y == 618) || (x == 523 && y == 7'd539) || (x == 7'd5 && y == 7'd151) ||
		(x == 7'd410 && y == 7'd175) || (x == 291 && y == 155) || (x == 347 && y == 7'd348) ||
		(x == 7'd42 && y == 550) || (x == 70 && y == 7) || (x == 7'd617 && y == 7'd112) ||
		(x == 369 && y == 632) || (x == 7'd304 && y == 7'd131) || (x == 636 && y == 7'd172) ||
		(x == 7'd561 && y == 7'd144) || (x == 7'd334 && y == 7'd603) || (x == 7'd417 && y == 86) ||
		(x == 184 && y == 302) || (x == 7'd171 && y == 7'd595) || (x == 493 && y == 7'd372) ||
		(x == 7'd569 && y == 7'd194) || (x == 104 && y == 7'd331) || (x == 245 && y == 192) ||
		(x == 7'd38 && y == 182) || (x == 7'd316 && y == 205) || (x == 7'd371 && y == 7'd313) ||
		(x == 7'd419 && y == 7'd346) || (x == 242 && y == 545) || (x == 7'd117 && y == 479) ||
		(x == 380 && y == 7'd36) || (x == 7'd571 && y == 7'd198) || (x == 7'd560 && y == 7'd394) ||
		(x == 7'd229 && y == 7'd553) || (x == 7'd208 && y == 7'd497) || (x == 7'd474 && y == 7'd337) ||
		(x == 7'd6 && y == 592) || (x == 7'd266 && y == 7'd569) || (x == 7'd356 && y == 7'd298) ||
		(x == 7'd217 && y == 7'd377) || (x == 7'd244 && y == 7'd198) || (x == 7'd615 && y == 602) ||
		(x == 565 && y == 179) || (x == 417 && y == 7'd382) || (x == 200 && y == 7'd356) ||
		(x == 7'd456 && y == 15) || (x == 576 && y == 7'd53) || (x == 7'd63 && y == 7'd211) ||
		(x == 7'd125 && y == 25) || (x == 7'd4 && y == 7'd606) || (x == 518 && y == 518) ||
		(x == 7'd590 && y == 298) || (x == 602 && y == 399) || (x == 446 && y == 452) ||
		(x == 7'd153 && y == 7'd523) || (x == 496 && y == 7'd492) || (x == 401 && y == 7'd274) ||
		(x == 516 && y == 311) || (x == 457 && y == 385) || (x == 342 && y == 7'd364) ||
		(x == 484 && y == 7'd154) || (x == 460 && y == 376) || (x == 7'd326 && y == 7'd546) ||
		(x == 7'd190 && y == 7'd611) || (x == 481 && y == 197) || (x == 7'd104 && y == 7'd611) ||
		(x == 490 && y == 371) || (x == 7'd296 && y == 321) || (x == 159 && y == 466) ||
		(x == 445 && y == 7'd161) || (x == 350 && y == 7'd361) || (x == 7'd551 && y == 7'd391) ||
		(x == 7'd571 && y == 7'd323) || (x == 7'd269 && y == 64) || (x == 327 && y == 7'd207) ||
		(x == 153 && y == 557) || (x == 7'd527 && y == 589) || (x == 7'd151 && y == 7'd414) ||
		(x == 309 && y == 7'd146) || (x == 7'd52 && y == 153) || (x == 531 && y == 7'd188) ||
		(x == 7'd17 && y == 570) || (x == 185 && y == 294) || (x == 7'd190 && y == 619) ||
		(x == 224 && y == 396) || (x == 220 && y == 433) || (x == 7'd15 && y == 7'd530) ||
		(x == 150 && y == 252) || (x == 7'd144 && y == 7'd469) || (x == 329 && y == 7'd528) ||
		(x == 7'd535 && y == 402) || (x == 7'd404 && y == 263) || (x == 168 && y == 7'd332) ||
		(x == 7'd327 && y == 242) || (x == 546 && y == 7'd483) || (x == 565 && y == 7'd321) ||
		(x == 121 && y == 7'd142) || (x == 7'd573 && y == 7'd140) || (x == 7'd158 && y == 501) ||
		(x == 7'd583 && y == 477) || (x == 7'd326 && y == 248) || (x == 7'd565 && y == 25) ||
		(x == 7'd318 && y == 285) || (x == 7'd579 && y == 7'd40) || (x == 7'd42 && y == 312) ||
		(x == 476 && y == 538) || (x == 7'd576 && y == 376) || (x == 381 && y == 303) ||
		(x == 155 && y == 290) || (x == 562 && y == 440) || (x == 7'd406 && y == 7'd390) ||
		(x == 7'd37 && y == 287) || (x == 476 && y == 7'd9) || (x == 7'd210 && y == 7'd156) ||
		(x == 7'd229 && y == 7'd16) || (x == 7'd627 && y == 7'd238) || (x == 7'd502 && y == 7'd456) ||
		(x == 7'd4 && y == 270) || (x == 7'd180 && y == 375) || (x == 253 && y == 7'd527) ||
		(x == 7'd517 && y == 7'd451) || (x == 7'd570 && y == 7'd216) || (x == 320 && y == 7'd562) ||
		(x == 7'd276 && y == 7'd176) || (x == 382 && y == 7'd540) || (x == 7'd181 && y == 512) ||
		(x == 7'd381 && y == 7'd535) || (x == 371 && y == 292) || (x == 7'd552 && y == 7'd397) ||
		(x == 473 && y == 7'd51) || (x == 7'd617 && y == 7'd213) || (x == 259 && y == 288) ||
		(x == 371 && y == 373) || (x == 7'd47 && y == 487) || (x == 7'd251 && y == 436) ||
		(x == 292 && y == 415) || (x == 7'd362 && y == 304) || (x == 7'd502 && y == 7'd269) ||
		(x == 7'd353 && y == 323) || (x == 7'd218 && y == 7'd507) || (x == 320 && y == 434) ||
		(x == 7'd609 && y == 7'd294) || (x == 7'd454 && y == 7'd617) || (x == 312 && y == 424) ||
		(x == 7'd524 && y == 61) || (x == 626 && y == 7'd213) || (x == 7'd346 && y == 7'd346) ||
		(x == 196 && y == 441) || (x == 7'd511 && y == 216) || (x == 7'd338 && y == 7'd249) ||
		(x == 370 && y == 7'd582) || (x == 607 && y == 533) || (x == 7'd527 && y == 83) ||
		(x == 462 && y == 7'd93) || (x == 502 && y == 318) || (x == 7'd458 && y == 396) ||
		(x == 254 && y == 562) || (x == 417 && y == 536) || (x == 470 && y == 340) ||
		(x == 556 && y == 7'd310) || (x == 7'd508 && y == 7'd250) || (x == 174 && y == 7'd8) ||
		(x == 7'd637 && y == 7'd595) || (x == 554 && y == 238) || (x == 203 && y == 385) ||
		(x == 7'd423 && y == 7'd395) || (x == 7'd363 && y == 553) || (x == 7'd528 && y == 7'd385) ||
		(x == 478 && y == 7'd278) || (x == 7'd98 && y == 395) || (x == 569 && y == 7'd219) ||
		(x == 522 && y == 179) || (x == 7'd243 && y == 12) || (x == 7'd318 && y == 7'd140) ||
		(x == 7'd450 && y == 162) || (x == 7'd132 && y == 265) || (x == 109 && y == 7'd424) ||
		(x == 7'd459 && y == 7'd470) || (x == 447 && y == 7'd518) || (x == 411 && y == 197) ||
		(x == 7'd178 && y == 7'd385) || (x == 443 && y == 163) || (x == 7'd242 && y == 7'd29) ||
		(x == 7'd474 && y == 7'd133) || (x == 275 && y == 7'd235) || (x == 225 && y == 352) ||
		(x == 584 && y == 7'd368) || (x == 7'd554 && y == 7'd494) || (x == 7'd225 && y == 40) ||
		(x == 453 && y == 581) || (x == 7'd243 && y == 230) || (x == 7'd398 && y == 7'd496) ||
		(x == 7'd343 && y == 444) || (x == 326 && y == 7'd423) || (x == 7'd286 && y == 7'd72) ||
		(x == 7'd354 && y == 7'd530) || (x == 480 && y == 7'd369) || (x == 469 && y == 515) ||
		(x == 468 && y == 7'd573) || (x == 454 && y == 531) || (x == 7'd337 && y == 429) ||
		(x == 7'd160 && y == 386) || (x == 7'd453 && y == 7'd124) || (x == 20 && y == 77) ||
		(x == 7'd223 && y == 7'd544) || (x == 7'd283 && y == 7'd39) || (x == 7'd362 && y == 225) ||
		(x == 7'd594 && y == 360) || (x == 7'd81 && y == 575) || (x == 7'd490 && y == 132) ||
		(x == 317 && y == 7'd3) || (x == 7'd4 && y == 7'd391) || (x == 7'd540 && y == 151) ||
		(x == 7'd113 && y == 7'd494) || (x == 7'd15 && y == 7'd38) || (x == 7'd553 && y == 605) ||
		(x == 7'd424 && y == 7'd371) || (x == 363 && y == 7'd639) || (x == 7'd390 && y == 149) ||
		(x == 7'd103 && y == 360) || (x == 314 && y == 7'd428) || (x == 7'd144 && y == 7'd386) ||
		(x == 214 && y == 7'd305) || (x == 407 && y == 402) || (x == 485 && y == 7'd271) ||
		(x == 7'd220 && y == 29) || (x == 65 && y == 7'd609) || (x == 7'd519 && y == 7'd302) ||
		(x == 157 && y == 572) || (x == 314 && y == 7'd183) || (x == 7'd362 && y == 49) ||
		(x == 7'd141 && y == 7'd17) || (x == 7'd342 && y == 7'd628) || (x == 7'd283 && y == 7'd635) ||
		(x == 404 && y == 7'd419) || (x == 429 && y == 7'd277) || (x == 3 && y == 7'd457) ||
		(x == 7'd524 && y == 467) || (x == 304 && y == 136) || (x == 196 && y == 143) ||
		(x == 7'd398 && y == 492) || (x == 571 && y == 569) || (x == 164 && y == 7'd622) ||
		(x == 7'd156 && y == 7'd44) || (x == 138 && y == 462) || (x == 7'd351 && y == 158) ||
		(x == 7'd452 && y == 7'd508) || (x == 7'd321 && y == 7'd605) || (x == 450 && y == 7'd307) ||
		(x == 7'd344 && y == 7'd284) || (x == 7'd611 && y == 55) || (x == 321 && y == 211) ||
		(x == 7'd523 && y == 420) || (x == 633 && y == 484) || (x == 281 && y == 7'd126) ||
		(x == 7'd561 && y == 125) || (x == 191 && y == 7'd501) || (x == 127 && y == 7'd387) ||
		(x == 7'd625 && y == 7'd273) || (x == 130 && y == 7'd126) || (x == 188 && y == 7'd251) ||
		(x == 204 && y == 172) || (x == 7'd125 && y == 7'd404) || (x == 307 && y == 286) ||
		(x == 7'd618 && y == 521) || (x == 7'd222 && y == 7'd420) || (x == 27 && y == 7'd125) ||
		(x == 7'd535 && y == 7'd437) || (x == 423 && y == 526) || (x == 7'd602 && y == 7'd485) ||
		(x == 304 && y == 7'd318) || (x == 536 && y == 7'd502) || (x == 7'd486 && y == 337) ||
		(x == 7'd410 && y == 7'd408) || (x == 7'd522 && y == 7'd575) || (x == 536 && y == 7'd567) ||
		(x == 282 && y == 7'd551) || (x == 7'd9 && y == 516) || (x == 230 && y == 326) ||
		(x == 7'd548 && y == 7'd241) || (x == 7'd133 && y == 625) || (x == 7'd383 && y == 7'd115) ||
		(x == 7'd24 && y == 372) || (x == 499 && y == 7'd11) || (x == 294 && y == 194) ||
		(x == 142 && y == 151) || (x == 601 && y == 7'd605) || (x == 7'd603 && y == 7'd545) ||
		(x == 7'd595 && y == 7'd241) || (x == 114 && y == 7'd545) || (x == 169 && y == 7'd446) ||
		(x == 448 && y == 7'd369) || (x == 72 && y == 7'd591) || (x == 7'd553 && y == 224) ||
		(x == 7'd382 && y == 120) || (x == 509 && y == 7'd246) || (x == 171 && y == 532) ||
		(x == 581 && y == 7'd93) || (x == 520 && y == 7'd189) || (x == 475 && y == 7'd496) ||
		(x == 7'd621 && y == 583) || (x == 169 && y == 7'd443) || (x == 7'd68 && y == 7'd627) ||
		(x == 137 && y == 7'd568) || (x == 7'd145 && y == 7'd313) || (x == 7'd142 && y == 7'd501) ||
		(x == 7'd531 && y == 7'd133) || (x == 7'd517 && y == 7'd131) || (x == 7'd322 && y == 7'd79) ||
		(x == 7'd634 && y == 238) || (x == 7'd583 && y == 7'd527) || (x == 326 && y == 390) ||
		(x == 282 && y == 375) || (x == 7'd36 && y == 7'd118) || (x == 7'd150 && y == 7'd334) ||
		(x == 7'd82 && y == 493) || (x == 634 && y == 7'd226) || (x == 102 && y == 7'd369) ||
		(x == 267 && y == 7'd530) || (x == 7'd621 && y == 7'd599) || (x == 172 && y == 7'd213) ||
		(x == 192 && y == 7'd333) || (x == 508 && y == 363) || (x == 7'd510 && y == 7'd259) ||
		(x == 7'd388 && y == 7'd588) || (x == 262 && y == 226) || (x == 62 && y == 7'd500) ||
		(x == 7'd134 && y == 7'd279) || (x == 7'd502 && y == 407) || (x == 7'd130 && y == 298) ||
		(x == 7'd627 && y == 123) || (x == 7'd84 && y == 7'd499) || (x == 232 && y == 7'd155) ||
		(x == 7'd338 && y == 7'd380) || (x == 594 && y == 147) || (x == 350 && y == 546) ||
		(x == 7'd480 && y == 7'd466) || (x == 7'd377 && y == 201) || (x == 306 && y == 7'd236) ||
		(x == 581 && y == 242) || (x == 268 && y == 7'd343) || (x == 226 && y == 246) ||
		(x == 284 && y == 294) || (x == 7'd235 && y == 25) || (x == 261 && y == 581) ||
		(x == 7'd185 && y == 7'd90) || (x == 254 && y == 7'd282) || (x == 619 && y == 7'd589) ||
		(x == 7'd134 && y == 186) || (x == 7'd349 && y == 7'd600) || (x == 188 && y == 7'd555) ||
		(x == 7'd317 && y == 574) || (x == 7'd105 && y == 7'd613) || (x == 554 && y == 434) ||
		(x == 258 && y == 7'd494) || (x == 330 && y == 396) || (x == 7'd359 && y == 7'd539) ||
		(x == 7'd400 && y == 7'd131) || (x == 7'd468 && y == 7'd498) || (x == 412 && y == 538) ||
		(x == 7'd603 && y == 115) || (x == 607 && y == 7'd274) || (x == 123 && y == 7'd591) ||
		(x == 7'd114 && y == 7'd496) || (x == 140 && y == 440) || (x == 180 && y == 260) ||
		(x == 7'd203 && y == 7'd552) || (x == 7'd486 && y == 515) || (x == 321 && y == 7'd636) ||
		(x == 7'd4 && y == 596) || (x == 7'd138 && y == 64) || (x == 182 && y == 7'd28) ||
		(x == 182 && y == 519) || (x == 262 && y == 441) || (x == 7'd193 && y == 7'd584) ||
		(x == 7'd547 && y == 7'd447) || (x == 224 && y == 7'd631) || (x == 7'd304 && y == 7'd143) ||
		(x == 189 && y == 169) || (x == 7'd611 && y == 308) || (x == 73 && y == 7'd184) ||
		(x == 7'd344 && y == 344) || (x == 445 && y == 413) || (x == 520 && y == 515) ||
		(x == 518 && y == 441) || (x == 7'd120 && y == 7'd615) || (x == 111 && y == 7'd448) ||
		(x == 7'd520 && y == 408) || (x == 326 && y == 146) || (x == 578 && y == 7'd453) ||
		(x == 597 && y == 7'd614) || (x == 7'd65 && y == 7'd506) || (x == 7'd263 && y == 7'd196) ||
		(x == 182 && y == 394) || (x == 7'd177 && y == 577) || (x == 41 && y == 7'd181) ||
		(x == 161 && y == 314) || (x == 7'd312 && y == 7'd582) || (x == 484 && y == 255) ||
		(x == 434 && y == 607) || (x == 283 && y == 7'd455) || (x == 7'd367 && y == 7'd251) ||
		(x == 458 && y == 295) || (x == 623 && y == 617) || (x == 7'd259 && y == 101) ||
		(x == 7'd332 && y == 487) || (x == 7'd439 && y == 182) || (x == 445 && y == 7'd507) ||
		(x == 637 && y == 202) || (x == 7'd198 && y == 378) || (x == 401 && y == 7'd48) ||
		(x == 189 && y == 7'd625) || (x == 583 && y == 340) || (x == 7'd462 && y == 7'd251) ||
		(x == 326 && y == 529) || (x == 7'd410 && y == 7'd183) || (x == 451 && y == 182) ||
		(x == 7'd357 && y == 447) || (x == 7'd247 && y == 7'd353) || (x == 300 && y == 498) ||
		(x == 7'd163 && y == 7'd273) || (x == 7'd316 && y == 120) || (x == 334 && y == 7'd134) ||
		(x == 7'd506 && y == 7'd181) || (x == 283 && y == 584) || (x == 7'd243 && y == 7'd352) ||
		(x == 436 && y == 7'd270) || (x == 148 && y == 7'd131) || (x == 7'd307 && y == 7'd15) ||
		(x == 7'd277 && y == 586) || (x == 218 && y == 7'd607) || (x == 7'd401 && y == 7'd443) ||
		(x == 7'd498 && y == 120) || (x == 519 && y == 7'd301) || (x == 7'd521 && y == 7'd444) ||
		(x == 7'd615 && y == 7'd280) || (x == 7'd553 && y == 156) || (x == 167 && y == 443) ||
		(x == 7'd531 && y == 538) || (x == 7'd196 && y == 368) || (x == 164 && y == 7'd46) ||
		(x == 7'd539 && y == 7'd385) || (x == 7'd545 && y == 617) || (x == 7'd578 && y == 199) ||
		(x == 7'd583 && y == 7'd363) || (x == 7'd567 && y == 254) || (x == 7'd266 && y == 371) ||
		(x == 200 && y == 181) || (x == 7'd586 && y == 153) || (x == 221 && y == 7'd214) ||
		(x == 7'd459 && y == 43) || (x == 379 && y == 7'd200) || (x == 7'd602 && y == 7'd504) ||
		(x == 7'd97 && y == 384) || (x == 580 && y == 348) || (x == 365 && y == 7'd235) ||
		(x == 586 && y == 7'd115) || (x == 7'd148 && y == 313) || (x == 244 && y == 7'd109) ||
		(x == 480 && y == 7'd562) || (x == 252 && y == 186) || (x == 285 && y == 417) ||
		(x == 7'd516 && y == 420) || (x == 7'd16 && y == 165) || (x == 633 && y == 221) ||
		(x == 7'd184 && y == 422) || (x == 400 && y == 452) || (x == 234 && y == 7'd275) ||
		(x == 7'd391 && y == 7'd389) || (x == 335 && y == 7'd217) || (x == 7'd82 && y == 188) ||
		(x == 135 && y == 427) || (x == 603 && y == 224) || (x == 7'd8 && y == 167) ||
		(x == 310 && y == 7'd329) || (x == 160 && y == 7'd349) || (x == 7'd144 && y == 21) ||
		(x == 400 && y == 323) || (x == 412 && y == 7'd89) || (x == 7'd519 && y == 7'd256) ||
		(x == 240 && y == 579) || (x == 7'd560 && y == 7'd479) || (x == 7'd195 && y == 7'd184) ||
		(x == 7'd194 && y == 7'd371) || (x == 585 && y == 7'd275) || (x == 7'd262 && y == 7'd569) ||
		(x == 7'd361 && y == 7'd455) || (x == 7'd279 && y == 7'd176) || (x == 7'd335 && y == 7'd508) ||
		(x == 7'd178 && y == 397) || (x == 7'd367 && y == 93) || (x == 7'd71 && y == 7'd436) ||
		(x == 7'd559 && y == 7'd133) || (x == 110 && y == 7'd180) || (x == 7'd196 && y == 7'd334) ||
		(x == 7'd620 && y == 7'd258) || (x == 7'd198 && y == 383) || (x == 7'd170 && y == 7'd284) ||
		(x == 7'd201 && y == 7'd146) || (x == 568 && y == 339) || (x == 7'd381 && y == 7'd514) ||
		(x == 7'd371 && y == 7'd414) || (x == 386 && y == 7'd634) || (x == 415 && y == 7'd54) ||
		(x == 7'd624 && y == 202) || (x == 58 && y == 7'd610) || (x == 7'd598 && y == 471) ||
		(x == 7'd130 && y == 7'd483) || (x == 7'd288 && y == 7'd19) || (x == 607 && y == 174) ||
		(x == 270 && y == 210) || (x == 454 && y == 247) || (x == 318 && y == 331) ||
		(x == 7'd633 && y == 246) || (x == 7'd517 && y == 7'd159) || (x == 492 && y == 7'd609) ||
		(x == 212 && y == 7'd535) || (x == 7'd372 && y == 7'd237) || (x == 7'd563 && y == 154) ||
		(x == 387 && y == 7'd456) || (x == 7'd14 && y == 7'd39) || (x == 7'd429 && y == 348) ||
		(x == 7'd390 && y == 3) || (x == 7'd248 && y == 7'd470) || (x == 7'd30 && y == 7'd515) ||
		(x == 194 && y == 7'd280) || (x == 507 && y == 244) || (x == 639 && y == 447) ||
		(x == 68 && y == 7'd177) || (x == 322 && y == 399) || (x == 624 && y == 444) ||
		(x == 223 && y == 7'd14) || (x == 7'd229 && y == 7'd332) || (x == 7'd112 && y == 592) ||
		(x == 399 && y == 424) || (x == 270 && y == 612) || (x == 566 && y == 222) ||
		(x == 60 && y == 7'd399) || (x == 487 && y == 7'd27) || (x == 7'd138 && y == 7'd169) ||
		(x == 7'd466 && y == 418) || (x == 7'd85 && y == 7'd427) || (x == 328 && y == 450) ||
		(x == 620 && y == 7'd398) || (x == 7'd435 && y == 144) || (x == 7'd278 && y == 7'd435) ||
		(x == 316 && y == 7'd547) || (x == 504 && y == 7'd483) || (x == 7'd472 && y == 7'd136) ||
		(x == 7'd221 && y == 232) || (x == 547 && y == 386) || (x == 7'd344 && y == 539) ||
		(x == 64 && y == 7'd560) || (x == 574 && y == 357) || (x == 7'd594 && y == 7'd358) ||
		(x == 7'd631 && y == 7'd226) || (x == 555 && y == 7'd231) || (x == 7'd526 && y == 7'd216) ||
		(x == 7'd579 && y == 490) || (x == 7'd530 && y == 7'd400) || (x == 503 && y == 7'd197) ||
		(x == 387 && y == 272) || (x == 7'd234 && y == 347) || (x == 493 && y == 567) ||
		(x == 7'd70 && y == 137) || (x == 7'd170 && y == 7'd239) || (x == 7'd502 && y == 7'd417) ||
		(x == 153 && y == 7'd173) || (x == 7'd200 && y == 7'd549) || (x == 7'd441 && y == 7'd239) ||
		(x == 147 && y == 271) || (x == 7'd440 && y == 7'd509) || (x == 495 && y == 622) ||
		(x == 115 && y == 7'd159) || (x == 492 && y == 7'd103) || (x == 330 && y == 7'd320) ||
		(x == 7'd389 && y == 7'd569) || (x == 200 && y == 610) || (x == 7'd529 && y == 7'd375) ||
		(x == 7'd314 && y == 7'd258) || (x == 406 && y == 7'd363) || (x == 145 && y == 237) ||
		(x == 148 && y == 7'd455) || (x == 508 && y == 341) || (x == 144 && y == 7'd162) ||
		(x == 629 && y == 203) || (x == 7'd621 && y == 7'd351) || (x == 7'd366 && y == 327) ||
		(x == 7'd145 && y == 33) || (x == 7'd521 && y == 439) || (x == 537 && y == 195) ||
		(x == 7'd356 && y == 110) || (x == 308 && y == 7'd500) || (x == 7'd405 && y == 7'd300) ||
		(x == 390 && y == 165) || (x == 7'd402 && y == 7'd494) || (x == 7'd274 && y == 7'd632) ||
		(x == 432 && y == 7'd353) || (x == 7'd407 && y == 345) || (x == 7'd422 && y == 7'd341) ||
		(x == 7'd146 && y == 7'd496) || (x == 255 && y == 7'd92) || (x == 475 && y == 7'd159) ||
		(x == 7'd615 && y == 7'd487) || (x == 7'd379 && y == 236) || (x == 257 && y == 7'd630) ||
		(x == 197 && y == 256) || (x == 407 && y == 7'd280) || (x == 7'd590 && y == 213) ||
		(x == 7'd347 && y == 506) || (x == 7'd466 && y == 7'd47) || (x == 7'd131 && y == 7'd196) ||
		(x == 7'd134 && y == 7'd134) || (x == 7'd177 && y == 237) || (x == 256 && y == 7'd577) ||
		(x == 7'd578 && y == 303) || (x == 470 && y == 396) || (x == 591 && y == 7'd237) ||
		(x == 207 && y == 7'd545) || (x == 7'd463 && y == 449) || (x == 7'd277 && y == 7'd466) ||
		(x == 576 && y == 212) || (x == 7'd334 && y == 7'd542) || (x == 7'd199 && y == 254) ||
		(x == 7'd616 && y == 7'd514) || (x == 7'd321 && y == 453) || (x == 210 && y == 7'd102) ||
		(x == 7'd342 && y == 7'd85) || (x == 7'd411 && y == 7'd438) || (x == 7'd468 && y == 264) ||
		(x == 7'd234 && y == 7'd470) || (x == 7'd290 && y == 7'd220) || (x == 277 && y == 7'd567) ||
		(x == 7'd107 && y == 7'd497) || (x == 309 && y == 413) || (x == 25 && y == 7'd617) ||
		(x == 26 && y == 7'd178) || (x == 7'd369 && y == 7'd91) || (x == 64 && y == 91) ||
		(x == 21 && y == 7'd158) || (x == 7'd321 && y == 7'd324) || (x == 7'd127 && y == 241) ||
		(x == 541 && y == 227) || (x == 7'd317 && y == 569) || (x == 97 && y == 7'd523) ||
		(x == 7'd259 && y == 7'd565) || (x == 7'd117 && y == 7'd519) || (x == 7'd376 && y == 7'd316) ||
		(x == 622 && y == 7'd81) || (x == 493 && y == 436) || (x == 7'd434 && y == 7'd550) ||
		(x == 7'd613 && y == 7'd465) || (x == 319 && y == 7'd34) || (x == 7'd484 && y == 7'd532) ||
		(x == 142 && y == 466) || (x == 7'd338 && y == 265) || (x == 7'd449 && y == 37) ||
		(x == 450 && y == 7'd378) || (x == 7'd248 && y == 7'd412) || (x == 7'd73 && y == 2) ||
		(x == 7'd154 && y == 7'd10) || (x == 275 && y == 7'd596) || (x == 7'd245 && y == 309) ||
		(x == 7'd370 && y == 7'd6) || (x == 7'd146 && y == 7'd566) || (x == 7'd308 && y == 7'd355) ||
		(x == 182 && y == 519) || (x == 365 && y == 7'd574) || (x == 7'd633 && y == 7'd550) ||
		(x == 68 && y == 7'd309) || (x == 292 && y == 7'd633) || (x == 280 && y == 7'd134) ||
		(x == 277 && y == 624) || (x == 7'd542 && y == 7'd396) || (x == 7'd498 && y == 7'd310) ||
		(x == 7'd616 && y == 7'd340) || (x == 7'd133 && y == 393) || (x == 7'd585 && y == 459) ||
		(x == 166 && y == 7'd163) || (x == 7'd423 && y == 7'd625) || (x == 356 && y == 7'd319) ||
		(x == 292 && y == 197) || (x == 357 && y == 7'd231) || (x == 7'd413 && y == 227) ||
		(x == 7'd416 && y == 7'd505) || (x == 292 && y == 267) || (x == 7'd350 && y == 264) ||
		(x == 7'd231 && y == 7'd110) || (x == 7'd373 && y == 7'd35) || (x == 244 && y == 7'd191) ||
		(x == 7'd632 && y == 470) || (x == 7'd495 && y == 7'd515) || (x == 24 && y == 7'd135) ||
		(x == 475 && y == 553) || (x == 393 && y == 390) || (x == 296 && y == 7'd223) ||
		(x == 7'd454 && y == 7'd395) || (x == 540 && y == 7'd5) || (x == 7'd565 && y == 7'd528) ||
		(x == 146 && y == 206) || (x == 561 && y == 7'd379) || (x == 7'd181 && y == 7'd515) ||
		(x == 7'd367 && y == 7'd38) || (x == 7'd83 && y == 7'd50) || (x == 49 && y == 7'd382) ||
		(x == 7'd285 && y == 105) || (x == 7'd324 && y == 273) || (x == 7'd393 && y == 7'd473) ||
		(x == 7'd319 && y == 7'd504) || (x == 382 && y == 193) || (x == 435 && y == 7'd8) ||
		(x == 404 && y == 575) || (x == 382 && y == 509) || (x == 7'd80 && y == 7'd512) ||
		(x == 477 && y == 7'd543) || (x == 7'd152 && y == 7'd139) || (x == 159 && y == 576) ||
		(x == 503 && y == 7'd216) || (x == 184 && y == 7'd359) || (x == 487 && y == 7'd142) ||
		(x == 367 && y == 236) || (x == 132 && y == 414) || (x == 43 && y == 7'd637) ||
		(x == 241 && y == 237) || (x == 7'd277 && y == 7'd561) || (x == 7'd182 && y == 522) ||
		(x == 7'd593 && y == 7'd367) || (x == 7'd315 && y == 7'd531) || (x == 458 && y == 7'd482) ||
		(x == 7'd205 && y == 7'd366) || (x == 385 && y == 7'd575) || (x == 7'd362 && y == 7'd469) ||
		(x == 7'd501 && y == 7'd479) || (x == 259 && y == 7'd240) || (x == 219 && y == 521) ||
		(x == 7'd216 && y == 137) || (x == 307 && y == 7'd70) || (x == 413 && y == 372) ||
		(x == 311 && y == 277) || (x == 607 && y == 7'd535) || (x == 7'd366 && y == 7'd144) ||
		(x == 7'd240 && y == 7'd628) || (x == 7'd88 && y == 7'd4) || (x == 7'd84 && y == 590) ||
		(x == 7'd314 && y == 7'd369) || (x == 7'd148 && y == 7'd339) || (x == 7'd410 && y == 7'd222) ||
		(x == 532 && y == 7'd256) || (x == 277 && y == 291) || (x == 7'd409 && y == 7'd179) ||
		(x == 7'd459 && y == 7'd258) || (x == 7'd249 && y == 7'd568) || (x == 7'd448 && y == 404) ||
		(x == 209 && y == 7'd42) || (x == 7'd261 && y == 7'd249) || (x == 7'd383 && y == 7'd613) ||
		(x == 565 && y == 136) || (x == 7'd144 && y == 7'd13) || (x == 530 && y == 7'd612) ||
		(x == 7'd23 && y == 306) || (x == 7'd54 && y == 7'd286) || (x == 7'd599 && y == 7'd279) ||
		(x == 7'd477 && y == 632) || (x == 7'd337 && y == 320) || (x == 616 && y == 233) ||
		(x == 7'd196 && y == 113) || (x == 7'd373 && y == 7'd394) || (x == 478 && y == 7'd338) ||
		(x == 241 && y == 533) || (x == 442 && y == 7'd279) || (x == 531 && y == 7'd141) ||
		(x == 7'd514 && y == 7'd564) || (x == 7'd387 && y == 509) || (x == 409 && y == 332) ||
		(x == 143 && y == 567) || (x == 547 && y == 264) || (x == 7'd177 && y == 512) ||
		(x == 7'd499 && y == 226) || (x == 7'd537 && y == 290) || (x == 440 && y == 360) ||
		(x == 301 && y == 586) || (x == 270 && y == 536) || (x == 7'd346 && y == 7'd402) ||
		(x == 154 && y == 208) || (x == 7'd288 && y == 7'd592) || (x == 398 && y == 7'd384) ||
		(x == 7'd339 && y == 105) || (x == 381 && y == 7'd398) || (x == 376 && y == 7'd430) ||
		(x == 7'd355 && y == 7'd9) || (x == 7'd363 && y == 7'd601) || (x == 555 && y == 416) ||
		(x == 7'd577 && y == 7'd351) || (x == 593 && y == 7'd612) || (x == 7'd621 && y == 446) ||
		(x == 201 && y == 328) || (x == 7'd588 && y == 7'd513) || (x == 7'd471 && y == 257) ||
		(x == 7'd333 && y == 7'd257) || (x == 7'd453 && y == 7'd12) || (x == 7'd79 && y == 7'd455) ||
		(x == 7'd356 && y == 7'd568) || (x == 7'd476 && y == 7'd77) || (x == 580 && y == 7'd618) ||
		(x == 7'd15 && y == 7'd244) || (x == 331 && y == 7'd544) || (x == 7'd541 && y == 513) ||
		(x == 7'd20 && y == 7'd160) || (x == 269 && y == 7'd621) || (x == 7'd73 && y == 7'd478) ||
		(x == 93 && y == 7'd334) || (x == 510 && y == 204) || (x == 7'd606 && y == 7'd125) ||
		(x == 16 && y == 7'd182) || (x == 7'd401 && y == 315) || (x == 7'd455 && y == 7'd184) ||
		(x == 310 && y == 7'd416) || (x == 7'd639 && y == 7'd182) || (x == 142 && y == 7'd315) ||
		(x == 7'd87 && y == 90) || (x == 7'd545 && y == 7'd531) || (x == 7'd305 && y == 7'd292) ||
		(x == 7'd354 && y == 7'd554) || (x == 7'd124 && y == 7'd64) || (x == 7'd216 && y == 7'd407) ||
		(x == 7'd23 && y == 560) || (x == 186 && y == 7'd497) || (x == 7'd533 && y == 325) ||
		(x == 7'd308 && y == 7'd619) || (x == 7'd632 && y == 7'd140) || (x == 7'd125 && y == 7'd612) ||
		(x == 168 && y == 157) || (x == 7'd273 && y == 264) || (x == 7'd526 && y == 7'd402) ||
		(x == 562 && y == 386) || (x == 137 && y == 283) || (x == 573 && y == 7'd360) ||
		(x == 7'd184 && y == 262) || (x == 332 && y == 148) || (x == 7'd618 && y == 574) ||
		(x == 369 && y == 7'd610) || (x == 7'd154 && y == 7'd351) || (x == 7'd7 && y == 471) ||
		(x == 7'd110 && y == 451) || (x == 7'd311 && y == 185) || (x == 553 && y == 7'd139) ||
		(x == 115 && y == 7'd202) || (x == 7'd243 && y == 7'd478) || (x == 7'd317 && y == 7'd482) ||
		(x == 7'd97 && y == 338) || (x == 7'd481 && y == 181) || (x == 632 && y == 225) ||
		(x == 7'd166 && y == 7'd270) || (x == 196 && y == 7'd8) || (x == 421 && y == 7'd601) ||
		(x == 7'd91 && y == 291) || (x == 256 && y == 7'd104) || (x == 453 && y == 7'd166) ||
		(x == 225 && y == 274) || (x == 7'd598 && y == 7'd596) || (x == 628 && y == 7'd200) ||
		(x == 174 && y == 7'd60) || (x == 552 && y == 7'd224) || (x == 75 && y == 7'd298) ||
		(x == 337 && y == 428) || (x == 181 && y == 237) || (x == 7'd474 && y == 441) ||
		(x == 565 && y == 7'd423) || (x == 86 && y == 7'd389) || (x == 129 && y == 399) ||
		(x == 7'd382 && y == 66) || (x == 475 && y == 7'd100) || (x == 424 && y == 555) ||
		(x == 501 && y == 363) || (x == 7'd422 && y == 7'd3) || (x == 7'd464 && y == 7'd371) ||
		(x == 7'd422 && y == 114) || (x == 7'd358 && y == 7'd425) || (x == 495 && y == 7'd350) ||
		(x == 7'd82 && y == 87) || (x == 7'd86 && y == 102) || (x == 7'd543 && y == 13) ||
		(x == 60 && y == 7'd241) || (x == 549 && y == 302) || (x == 7'd626 && y == 7'd268) ||
		(x == 405 && y == 584) || (x == 7'd76 && y == 511) || (x == 480 && y == 7'd544) ||
		(x == 7'd382 && y == 7'd388) || (x == 7'd133 && y == 45) || (x == 201 && y == 399) ||
		(x == 7'd580 && y == 7'd562) || (x == 614 && y == 7'd297) || (x == 446 && y == 7'd192) ||
		(x == 460 && y == 348) || (x == 7'd469 && y == 7'd256) || (x == 7'd442 && y == 7'd276) ||
		(x == 7'd198 && y == 7'd417) || (x == 636 && y == 7'd317) || (x == 7'd26 && y == 7'd11) ||
		(x == 558 && y == 7'd399) || (x == 7'd504 && y == 7'd84) || (x == 325 && y == 7'd512) ||
		(x == 7'd173 && y == 235) || (x == 619 && y == 7'd440) || (x == 51 && y == 105) ||
		(x == 7'd334 && y == 7'd176) || (x == 7'd508 && y == 189) || (x == 7'd294 && y == 7'd529) ||
		(x == 511 && y == 7'd621) || (x == 443 && y == 7'd155) || (x == 7'd492 && y == 7'd606) ||
		(x == 7'd140 && y == 7'd466) || (x == 7'd251 && y == 242) || (x == 204 && y == 7'd448) ||
		(x == 7'd292 && y == 7'd144) || (x == 7'd104 && y == 193) || (x == 7'd583 && y == 7'd635) ||
		(x == 7'd165 && y == 372) || (x == 7'd332 && y == 7'd160) || (x == 7'd365 && y == 30) ||
		(x == 7'd77 && y == 152) || (x == 7'd508 && y == 7'd324) || (x == 7'd14 && y == 476) ||
		(x == 7'd64 && y == 7'd447) || (x == 7'd301 && y == 7'd633) || (x == 537 && y == 219) ||
		(x == 7'd480 && y == 125) || (x == 7'd453 && y == 7'd180) || (x == 7'd409 && y == 298) ||
		(x == 199 && y == 284) || (x == 7'd329 && y == 7'd52) || (x == 225 && y == 7'd386) ||
		(x == 7'd387 && y == 7'd564) || (x == 7'd24 && y == 302) || (x == 7'd131 && y == 7'd154) ||
		(x == 203 && y == 7'd33) || (x == 7'd403 && y == 7'd150) || (x == 559 && y == 145) ||
		(x == 7'd444 && y == 7'd448) || (x == 7'd517 && y == 7'd288) || (x == 351 && y == 577) ||
		(x == 245 && y == 437) || (x == 7'd572 && y == 591) || (x == 153 && y == 7'd25) ||
		(x == 507 && y == 7'd567) || (x == 7'd517 && y == 7'd142) || (x == 286 && y == 364) ||
		(x == 494 && y == 538) || (x == 463 && y == 7'd116) || (x == 7'd66 && y == 7'd173) ||
		(x == 7'd235 && y == 602) || (x == 409 && y == 7'd210) || (x == 313 && y == 425) ||
		(x == 7'd510 && y == 149) || (x == 391 && y == 7'd295) || (x == 7'd511 && y == 376) ||
		(x == 223 && y == 7'd38) || (x == 7'd141 && y == 7'd342) || (x == 7'd452 && y == 349) ||
		(x == 7'd415 && y == 433) || (x == 202 && y == 176) || (x == 7'd189 && y == 340) ||
		(x == 7'd325 && y == 151) || (x == 7'd179 && y == 520) || (x == 7'd177 && y == 388) ||
		(x == 7'd637 && y == 7'd274) || (x == 7'd597 && y == 7'd563) || (x == 7'd628 && y == 480) ||
		(x == 7'd233 && y == 7'd635) || (x == 7'd210 && y == 7'd449) || (x == 422 && y == 285) ||
		(x == 11 && y == 7'd348) || (x == 7'd338 && y == 455) || (x == 7'd421 && y == 295) ||
		(x == 7'd332 && y == 7'd553) || (x == 7'd477 && y == 393) || (x == 7'd271 && y == 509) ||
		(x == 7'd454 && y == 7'd525) || (x == 7'd382 && y == 83) || (x == 7'd470 && y == 561) ||
		(x == 410 && y == 309) || (x == 196 && y == 7'd274) || (x == 7'd271 && y == 7'd513) ||
		(x == 345 && y == 7'd6) || (x == 7'd426 && y == 7'd134) || (x == 512 && y == 398) ||
		(x == 213 && y == 468) || (x == 7'd126 && y == 7'd335) || (x == 7'd440 && y == 156) ||
		(x == 341 && y == 130) || (x == 59 && y == 7'd498) || (x == 7'd584 && y == 257) ||
		(x == 7'd105 && y == 7'd608) || (x == 7'd125 && y == 7'd147) || (x == 388 && y == 394) ||
		(x == 501 && y == 7'd338) || (x == 7'd120 && y == 425) || (x == 7'd466 && y == 7'd195) ||
		(x == 7'd21 && y == 7'd632) || (x == 7'd188 && y == 7'd450) || (x == 577 && y == 7'd208) ||
		(x == 7'd530 && y == 7'd397) || (x == 382 && y == 7'd599) || (x == 7'd264 && y == 7'd462) ||
		(x == 475 && y == 333) || (x == 7'd472 && y == 181) || (x == 7'd621 && y == 7'd260) ||
		(x == 553 && y == 7'd604) || (x == 290 && y == 7'd53) || (x == 7'd391 && y == 7'd329) ||
		(x == 100 && y == 7'd616) || (x == 579 && y == 574) || (x == 465 && y == 420) ||
		(x == 349 && y == 7'd451) || (x == 7'd118 && y == 7'd166) || (x == 596 && y == 7'd89) ||
		(x == 469 && y == 601) || (x == 381 && y == 565) || (x == 567 && y == 363) ||
		(x == 7'd336 && y == 7'd588) || (x == 340 && y == 7'd25) || (x == 91 && y == 7'd251) ||
		(x == 7'd341 && y == 7'd375) || (x == 7'd253 && y == 7'd360) || (x == 7'd595 && y == 7'd466) ||
		(x == 331 && y == 7'd6) || (x == 208 && y == 7'd323) || (x == 330 && y == 563) ||
		(x == 7'd348 && y == 394) || (x == 547 && y == 7'd513) || (x == 7'd53 && y == 452) ||
		(x == 7'd420 && y == 507) || (x == 522 && y == 395) || (x == 2 && y == 7'd614) ||
		(x == 253 && y == 7'd464) || (x == 7'd293 && y == 7'd548) || (x == 7'd95 && y == 558) ||
		(x == 417 && y == 462) || (x == 7'd543 && y == 518) || (x == 7'd305 && y == 416) ||
		(x == 361 && y == 286) || (x == 7'd357 && y == 7'd18) || (x == 7'd344 && y == 7'd424) ||
		(x == 135 && y == 7'd415) || (x == 7'd589 && y == 7'd175) || (x == 7'd214 && y == 7'd272) ||
		(x == 460 && y == 181) || (x == 293 && y == 540) || (x == 7'd365 && y == 7'd500) ||
		(x == 7'd34 && y == 446) || (x == 7'd194 && y == 7'd324) || (x == 395 && y == 410) ||
		(x == 7'd94 && y == 7'd207) || (x == 622 && y == 7'd135) || (x == 560 && y == 7'd34) ||
		(x == 7'd471 && y == 518) || (x == 7'd452 && y == 7'd189) || (x == 174 && y == 258) ||
		(x == 526 && y == 210) || (x == 7'd61 && y == 210) || (x == 7'd75 && y == 544) ||
		(x == 228 && y == 580) || (x == 7'd64 && y == 7'd449) || (x == 306 && y == 470) ||
		(x == 7'd105 && y == 7'd247) || (x == 7'd518 && y == 285) || (x == 470 && y == 7'd612) ||
		(x == 7'd76 && y == 389) || (x == 7'd328 && y == 148) || (x == 7'd443 && y == 29) ||
		(x == 507 && y == 7'd556) || (x == 7'd233 && y == 81) || (x == 479 && y == 7'd77) ||
		(x == 7'd330 && y == 437) || (x == 7'd627 && y == 7'd625) || (x == 164 && y == 218) ||
		(x == 7'd469 && y == 259) || (x == 529 && y == 7'd328) || (x == 7'd146 && y == 7'd440) ||
		(x == 437 && y == 311) || (x == 7'd165 && y == 7'd529) || (x == 559 && y == 340) ||
		(x == 449 && y == 175) || (x == 68 && y == 10) || (x == 7'd139 && y == 307) ||
		(x == 7'd345 && y == 36) || (x == 597 && y == 7'd553) || (x == 583 && y == 415) ||
		(x == 7'd388 && y == 7'd505) || (x == 7'd496 && y == 640) || (x == 7'd378 && y == 7'd294) ||
		(x == 7'd19 && y == 572) || (x == 7'd272 && y == 246) || (x == 7'd447 && y == 7'd15) ||
		(x == 232 && y == 7'd53) || (x == 7'd71 && y == 3) || (x == 219 && y == 7'd28) ||
		(x == 314 && y == 257) || (x == 7'd225 && y == 7'd419) || (x == 449 && y == 7'd128) ||
		(x == 595 && y == 7'd470) || (x == 7'd213 && y == 134) || (x == 7'd624 && y == 7'd218) ||
		(x == 7'd272 && y == 7'd595) || (x == 227 && y == 7'd335) || (x == 7'd262 && y == 7'd224) ||
		(x == 7'd157 && y == 7'd550) || (x == 148 && y == 296) || (x == 406 && y == 196) ||
		(x == 7'd293 && y == 157) || (x == 435 && y == 7'd281) || (x == 7'd13 && y == 364) ||
		(x == 571 && y == 7'd493) || (x == 7'd609 && y == 12) || (x == 517 && y == 7'd422) ||
		(x == 7'd507 && y == 7'd448) || (x == 570 && y == 499) || (x == 189 && y == 525) ||
		(x == 7'd559 && y == 7'd252) || (x == 7'd87 && y == 140) || (x == 7'd313 && y == 7'd252) ||
		(x == 7'd220 && y == 7'd249) || (x == 7'd52 && y == 615) || (x == 518 && y == 458) ||
		(x == 7'd233 && y == 7'd405) || (x == 7'd500 && y == 607) || (x == 7'd120 && y == 7'd313) ||
		(x == 7'd94 && y == 7'd394) || (x == 562 && y == 7'd522) || (x == 7'd152 && y == 428) ||
		(x == 381 && y == 491) || (x == 7'd366 && y == 7'd499) || (x == 206 && y == 7'd447) ||
		(x == 7'd558 && y == 293) || (x == 169 && y == 376) || (x == 569 && y == 542) ||
		(x == 521 && y == 7'd141) || (x == 7'd493 && y == 7'd349) || (x == 7'd485 && y == 7'd77) ||
		(x == 7'd462 && y == 7'd207) || (x == 7'd373 && y == 7'd421) || (x == 97 && y == 7'd232) ||
		(x == 58 && y == 7'd347) || (x == 350 && y == 209) || (x == 7'd594 && y == 7'd130) ||
		(x == 358 && y == 7'd153) || (x == 552 && y == 7'd599) || (x == 310 && y == 569) ||
		(x == 217 && y == 7'd14) || (x == 267 && y == 7'd135) || (x == 7'd240 && y == 7'd270) ||
		(x == 554 && y == 623) || (x == 7'd542 && y == 7'd208) || (x == 7'd484 && y == 141) ||
		(x == 611 && y == 520) || (x == 351 && y == 639) || (x == 560 && y == 235) ||
		(x == 7'd375 && y == 61) || (x == 7'd110 && y == 7'd27) || (x == 491 && y == 138) ||
		(x == 7'd10 && y == 7'd275) || (x == 7'd164 && y == 76) || (x == 7'd449 && y == 192) ||
		(x == 457 && y == 7'd288) || (x == 501 && y == 626) || (x == 328 && y == 457) ||
		(x == 364 && y == 7'd117) || (x == 7'd154 && y == 7'd261) || (x == 7'd24 && y == 506) ||
		(x == 7'd605 && y == 448) || (x == 7'd376 && y == 390) || (x == 7'd583 && y == 7'd513) ||
		(x == 290 && y == 286) || (x == 7'd418 && y == 7'd529) || (x == 7'd37 && y == 427) ||
		(x == 7'd536 && y == 238) || (x == 7'd500 && y == 216) || (x == 7'd196 && y == 7'd265) ||
		(x == 7'd300 && y == 7'd392) || (x == 142 && y == 7'd288) || (x == 7'd380 && y == 7'd210) ||
		(x == 7'd114 && y == 426) || (x == 520 && y == 152) || (x == 7'd637 && y == 256) ||
		(x == 310 && y == 7'd122) || (x == 256 && y == 303) || (x == 7'd89 && y == 7'd606) ||
		(x == 7'd400 && y == 7'd367) || (x == 241 && y == 302) || (x == 199 && y == 7'd11) ||
		(x == 7'd524 && y == 7'd548) || (x == 7'd407 && y == 80) || (x == 362 && y == 7'd417) ||
		(x == 625 && y == 476) || (x == 182 && y == 7'd588) || (x == 422 && y == 7'd625) ||
		(x == 265 && y == 7'd526) || (x == 124 && y == 7'd505) || (x == 7'd219 && y == 111) ||
		(x == 7'd91 && y == 605) || (x == 7'd556 && y == 202) || (x == 129 && y == 7'd514) ||
		(x == 368 && y == 443) || (x == 311 && y == 210) || (x == 192 && y == 7'd577) ||
		(x == 574 && y == 7'd73) || (x == 250 && y == 416) || (x == 162 && y == 340) ||
		(x == 7'd579 && y == 507) || (x == 7'd628 && y == 7'd184) || (x == 311 && y == 7'd403) ||
		(x == 154 && y == 7'd439) || (x == 251 && y == 551) || (x == 7'd638 && y == 226) ||
		(x == 553 && y == 7'd335) || (x == 629 && y == 7'd578) || (x == 599 && y == 214) ||
		(x == 7'd314 && y == 7'd345) || (x == 7'd539 && y == 355) || (x == 7'd64 && y == 152) ||
		(x == 7'd444 && y == 7'd556) || (x == 402 && y == 7'd457) || (x == 7'd394 && y == 7'd143) ||
		(x == 210 && y == 291) || (x == 405 && y == 7'd414) || (x == 7'd625 && y == 389) ||
		(x == 7'd357 && y == 7'd273) || (x == 7'd383 && y == 7'd375) || (x == 571 && y == 441) ||
		(x == 7'd135 && y == 7'd171) || (x == 7'd281 && y == 7'd8) || (x == 7'd445 && y == 7'd119) ||
		(x == 208 && y == 7'd579) || (x == 455 && y == 7'd487) || (x == 7'd187 && y == 7'd577) ||
		(x == 7'd436 && y == 7'd638) || (x == 562 && y == 7'd485) || (x == 108 && y == 7'd115) ||
		(x == 7'd181 && y == 7'd574) || (x == 7'd279 && y == 492) || (x == 7'd252 && y == 7'd613) ||
		(x == 292 && y == 514) || (x == 186 && y == 7'd447) || (x == 39 && y == 7'd388) ||
		(x == 7'd145 && y == 140) || (x == 253 && y == 452) || (x == 210 && y == 7'd470) ||
		(x == 7'd29 && y == 377) || (x == 7'd610 && y == 588) || (x == 7'd114 && y == 7'd224) ||
		(x == 17 && y == 7'd500) || (x == 7'd631 && y == 7'd585) || (x == 577 && y == 292) ||
		(x == 7'd631 && y == 7'd125) || (x == 7'd160 && y == 7'd163) || (x == 594 && y == 7'd433) ||
		(x == 7'd0 && y == 347) || (x == 428 && y == 7'd330) || (x == 7'd391 && y == 7'd323) ||
		(x == 7'd267 && y == 410) || (x == 7'd205 && y == 559) || (x == 254 && y == 141) ||
		(x == 137 && y == 620) || (x == 7'd192 && y == 7'd465) || (x == 7'd258 && y == 7'd229) ||
		(x == 555 && y == 472) || (x == 7'd247 && y == 7'd234) || (x == 7'd292 && y == 7'd617) ||
		(x == 487 && y == 7'd491) || (x == 7'd484 && y == 7'd624) || (x == 7'd134 && y == 7'd566) ||
		(x == 146 && y == 303) || (x == 7'd276 && y == 424) || (x == 7'd397 && y == 387) ||
		(x == 7'd122 && y == 229) || (x == 7'd129 && y == 178) || (x == 49 && y == 7'd233) ||
		(x == 7'd324 && y == 525) || (x == 7'd471 && y == 7'd345) || (x == 6 && y == 7'd222) ||
		(x == 436 && y == 7'd431) || (x == 552 && y == 7'd569) || (x == 7'd591 && y == 7'd431) ||
		(x == 563 && y == 7'd307) || (x == 511 && y == 7'd538) || (x == 7'd404 && y == 232) ||
		(x == 7'd334 && y == 112) || (x == 517 && y == 267) || (x == 419 && y == 7'd23) ||
		(x == 471 && y == 410) || (x == 7'd204 && y == 71) || (x == 7'd490 && y == 7'd426) ||
		(x == 432 && y == 288) || (x == 7'd17 && y == 7'd141) || (x == 7'd326 && y == 7'd464) ||
		(x == 7'd483 && y == 7'd614) || (x == 572 && y == 7'd522) || (x == 269 && y == 7'd270) ||
		(x == 7'd172 && y == 7'd635) || (x == 411 && y == 518) || (x == 356 && y == 7'd344) ||
		(x == 7'd397 && y == 333) || (x == 617 && y == 546) || (x == 78 && y == 7'd174) ||
		(x == 378 && y == 7'd493) || (x == 222 && y == 7'd514) || (x == 7'd453 && y == 7'd551) ||
		(x == 7'd193 && y == 7'd579) || (x == 7'd554 && y == 625) || (x == 7'd511 && y == 7'd299) ||
		(x == 276 && y == 7'd368) || (x == 342 && y == 245) || (x == 7'd272 && y == 7'd630) ||
		(x == 7'd620 && y == 7'd540) || (x == 7'd23 && y == 415) || (x == 485 && y == 288) ||
		(x == 505 && y == 7'd99) || (x == 7'd59 && y == 7'd347) || (x == 159 && y == 7'd535) ||
		(x == 634 && y == 188) || (x == 7'd388 && y == 7'd74) || (x == 7'd387 && y == 47) ||
		(x == 575 && y == 7'd43) || (x == 253 && y == 7'd310) || (x == 623 && y == 149) ||
		(x == 7'd19 && y == 632) || (x == 7'd210 && y == 497) || (x == 550 && y == 132) ||
		(x == 7'd216 && y == 7'd308) || (x == 157 && y == 7'd212) || (x == 191 && y == 7'd392) ||
		(x == 636 && y == 7'd45) || (x == 605 && y == 7'd299) || (x == 7'd440 && y == 550) ||
		(x == 479 && y == 598) || (x == 7'd399 && y == 7'd468) || (x == 278 && y == 7'd434) ||
		(x == 7'd411 && y == 582) || (x == 7'd327 && y == 7'd181) || (x == 7'd403 && y == 7'd629) ||
		(x == 67 && y == 90) || (x == 131 && y == 256) || (x == 7'd397 && y == 7'd245) ||
		(x == 502 && y == 7'd341) || (x == 57 && y == 7'd466) || (x == 603 && y == 179) ||
		(x == 291 && y == 391) || (x == 7'd519 && y == 7'd388) || (x == 7'd319 && y == 7'd553) ||
		(x == 7'd25 && y == 433) || (x == 7'd604 && y == 305) || (x == 7'd361 && y == 7'd278) ||
		(x == 394 && y == 628) || (x == 7'd590 && y == 631) || (x == 7'd410 && y == 101) ||
		(x == 7'd235 && y == 7'd298) || (x == 7'd452 && y == 604) || (x == 7'd267 && y == 155) ||
		(x == 232 && y == 605) || (x == 7'd532 && y == 278) || (x == 105 && y == 7'd371) ||
		(x == 7'd376 && y == 372) || (x == 438 && y == 306) || (x == 170 && y == 7'd201) ||
		(x == 7'd80 && y == 457) || (x == 7'd24 && y == 405) || (x == 7'd593 && y == 23) ||
		(x == 7'd442 && y == 7'd626) || (x == 7'd434 && y == 7'd274) || (x == 7'd629 && y == 426) ||
		(x == 7'd496 && y == 7'd477) || (x == 411 && y == 7'd392) || (x == 636 && y == 280) ||
		(x == 7'd212 && y == 7'd157) || (x == 7'd471 && y == 7'd604) || (x == 634 && y == 234) ||
		(x == 459 && y == 260) || (x == 167 && y == 7'd443) || (x == 7'd519 && y == 59) ||
		(x == 517 && y == 7'd582) || (x == 7'd224 && y == 7'd433) || (x == 7'd126 && y == 7'd182) ||
		(x == 7'd275 && y == 7'd377) || (x == 7'd164 && y == 7'd215) || (x == 7'd330 && y == 7'd131) ||
		(x == 308 && y == 7'd442) || (x == 406 && y == 633) || (x == 391 && y == 7'd578) ||
		(x == 7'd114 && y == 7'd627) || (x == 7'd7 && y == 400) || (x == 7'd32 && y == 7'd1) ||
		(x == 197 && y == 450) || (x == 575 && y == 269) || (x == 251 && y == 7'd219) ||
		(x == 210 && y == 460) || (x == 7'd319 && y == 395) || (x == 621 && y == 517) ||
		(x == 262 && y == 241) || (x == 543 && y == 7'd465) || (x == 489 && y == 7'd38) ||
		(x == 280 && y == 7'd432) || (x == 131 && y == 7'd190) || (x == 116 && y == 7'd183) ||
		(x == 7'd390 && y == 7'd395) || (x == 60 && y == 7'd388) || (x == 466 && y == 313) ||
		(x == 413 && y == 7'd539) || (x == 418 && y == 7'd416) || (x == 10 && y == 7'd632) ||
		(x == 65 && y == 7'd28) || (x == 240 && y == 546) || (x == 7'd73 && y == 233) ||
		(x == 304 && y == 344) || (x == 162 && y == 7'd284) || (x == 7'd501 && y == 611) ||
		(x == 7'd392 && y == 7'd473) || (x == 7'd383 && y == 7'd323) || (x == 7'd581 && y == 7'd131) ||
		(x == 485 && y == 331) || (x == 7'd64 && y == 7'd474) || (x == 269 && y == 619) ||
		(x == 7'd359 && y == 7'd336) || (x == 471 && y == 220) || (x == 7'd495 && y == 338) ||
		(x == 139 && y == 217) || (x == 7'd52 && y == 329) || (x == 7'd243 && y == 312) ||
		(x == 7'd238 && y == 7'd607) || (x == 7'd504 && y == 7'd573) || (x == 7'd25 && y == 181) ||
		(x == 7'd235 && y == 7'd44) || (x == 7'd350 && y == 519) || (x == 507 && y == 7'd623) ||
		(x == 286 && y == 621) || (x == 530 && y == 399) || (x == 7'd227 && y == 39) ||
		(x == 608 && y == 203) || (x == 638 && y == 7'd370) || (x == 466 && y == 7'd485) ||
		(x == 7'd276 && y == 70) || (x == 7'd622 && y == 89) || (x == 313 && y == 621) ||
		(x == 134 && y == 7'd162) || (x == 7'd470 && y == 71) || (x == 7'd568 && y == 323) ||
		(x == 7'd426 && y == 355) || (x == 404 && y == 7'd140) || (x == 7'd198 && y == 7'd591) ||
		(x == 7'd423 && y == 7'd134) || (x == 7'd53 && y == 551) || (x == 281 && y == 408) ||
		(x == 459 && y == 502) || (x == 7'd507 && y == 7'd449) || (x == 7'd612 && y == 7'd71) ||
		(x == 7'd273 && y == 7'd364) || (x == 7'd259 && y == 7'd438) || (x == 7'd60 && y == 7'd361) ||
		(x == 7'd398 && y == 483) || (x == 406 && y == 7'd108) || (x == 634 && y == 168) ||
		(x == 474 && y == 449) || (x == 261 && y == 7'd500) || (x == 418 && y == 7'd412) ||
		(x == 366 && y == 7'd48) || (x == 238 && y == 404) || (x == 265 && y == 7'd159) ||
		(x == 305 && y == 7'd401) || (x == 7'd525 && y == 268) || (x == 7'd263 && y == 7'd269) ||
		(x == 631 && y == 444) || (x == 488 && y == 129) || (x == 7'd316 && y == 262) ||
		(x == 7'd486 && y == 376) || (x == 7'd275 && y == 622) || (x == 7'd501 && y == 7'd264) ||
		(x == 7'd554 && y == 7'd617) || (x == 417 && y == 190) || (x == 7'd554 && y == 322) ||
		(x == 31 && y == 7'd453) || (x == 369 && y == 7'd234) || (x == 7'd105 && y == 173) ||
		(x == 7'd291 && y == 560) || (x == 7'd329 && y == 5) || (x == 7'd84 && y == 7'd363) ||
		(x == 575 && y == 357) || (x == 7'd326 && y == 7'd441) || (x == 7'd611 && y == 7'd275) ||
		(x == 450 && y == 131) || (x == 7'd623 && y == 114) || (x == 7'd244 && y == 319) ||
		(x == 7'd203 && y == 54) || (x == 7'd106 && y == 7'd24) || (x == 7'd548 && y == 247) ||
		(x == 132 && y == 179) || (x == 7'd209 && y == 414) || (x == 7'd290 && y == 91) ||
		(x == 7'd511 && y == 7'd536) || (x == 558 && y == 398) || (x == 7'd212 && y == 7'd583) ||
		(x == 430 && y == 7'd574) || (x == 163 && y == 7'd102) || (x == 7'd604 && y == 256) ||
		(x == 359 && y == 7'd405) || (x == 7'd503 && y == 7'd569) || (x == 264 && y == 549) ||
		(x == 328 && y == 7'd91) || (x == 7'd519 && y == 7'd416) || (x == 535 && y == 7'd521) ||
		(x == 518 && y == 7'd145) || (x == 7'd322 && y == 7'd245) || (x == 7'd486 && y == 7'd3) ||
		(x == 57 && y == 7'd491) || (x == 165 && y == 197) || (x == 7'd106 && y == 329) ||
		(x == 7'd369 && y == 221) || (x == 62 && y == 7'd318) || (x == 216 && y == 223) ||
		(x == 7'd254 && y == 7'd500) || (x == 331 && y == 7'd511) || (x == 7'd301 && y == 385) ||
		(x == 7'd137 && y == 161) || (x == 7'd469 && y == 554) || (x == 237 && y == 638) ||
		(x == 285 && y == 389) || (x == 431 && y == 534) || (x == 7'd438 && y == 7'd325) ||
		(x == 497 && y == 7'd69) || (x == 269 && y == 7'd156) || (x == 7'd274 && y == 485) ||
		(x == 7'd378 && y == 7'd446) || (x == 7'd508 && y == 504) || (x == 7'd321 && y == 328) ||
		(x == 278 && y == 281) || (x == 434 && y == 7'd255) || (x == 7'd110 && y == 7'd128) ||
		(x == 7'd573 && y == 7'd486) || (x == 7'd235 && y == 327) || (x == 7'd493 && y == 7'd299) ||
		(x == 7'd408 && y == 7'd392) || (x == 7'd488 && y == 584) || (x == 7'd393 && y == 7'd61) ||
		(x == 7'd558 && y == 39) || (x == 7'd397 && y == 497) || (x == 522 && y == 299) ||
		(x == 7'd329 && y == 7'd269) || (x == 186 && y == 569) || (x == 7'd386 && y == 31) ||
		(x == 7'd135 && y == 7'd386) || (x == 613 && y == 7'd389) || (x == 406 && y == 509) ||
		(x == 563 && y == 7'd197) || (x == 317 && y == 7'd329) || (x == 7'd141 && y == 7'd272) ||
		(x == 7'd400 && y == 562) || (x == 7'd39 && y == 577) || (x == 7'd489 && y == 7'd258) ||
		(x == 7'd341 && y == 7'd514) || (x == 268 && y == 7'd45) || (x == 7'd119 && y == 7'd136) ||
		(x == 7'd145 && y == 520) || (x == 588 && y == 145) || (x == 7'd402 && y == 0) ||
		(x == 7'd238 && y == 7'd181) || (x == 619 && y == 7'd61) || (x == 7'd355 && y == 7'd526) ||
		(x == 345 && y == 7'd33) || (x == 215 && y == 7'd188) || (x == 7'd148 && y == 7'd465) ||
		(x == 422 && y == 7'd593) || (x == 558 && y == 600) || (x == 298 && y == 7'd11) ||
		(x == 7'd5 && y == 145) || (x == 31 && y == 7'd557) || (x == 7'd436 && y == 7'd398) ||
		(x == 456 && y == 386) || (x == 518 && y == 227) || (x == 459 && y == 293) ||
		(x == 7'd497 && y == 194) || (x == 9 && y == 7'd443) || (x == 261 && y == 7'd151) ||
		(x == 7'd120 && y == 7'd460) || (x == 131 && y == 473) || (x == 7'd414 && y == 605) ||
		(x == 7'd168 && y == 7'd166) || (x == 158 && y == 7'd202) || (x == 7'd136 && y == 139) ||
		(x == 134 && y == 7'd127) || (x == 7'd371 && y == 7'd217) || (x == 21 && y == 7'd153) ||
		(x == 241 && y == 304) || (x == 319 && y == 7'd599) || (x == 7'd416 && y == 573) ||
		(x == 536 && y == 7'd240) || (x == 302 && y == 170) || (x == 176 && y == 494) ||
		(x == 7'd22 && y == 7'd394) || (x == 7'd410 && y == 530) || (x == 508 && y == 166) ||
		(x == 7'd206 && y == 7'd491) || (x == 7'd217 && y == 7'd469) || (x == 7'd73 && y == 7'd309) ||
		(x == 467 && y == 7'd65) || (x == 213 && y == 7'd213) || (x == 516 && y == 406) ||
		(x == 4 && y == 7'd395) || (x == 7'd50 && y == 7'd259) || (x == 345 && y == 7'd68) ||
		(x == 7'd299 && y == 7'd269) || (x == 7'd222 && y == 7'd215) || (x == 460 && y == 538) ||
		(x == 7'd9 && y == 591) || (x == 7'd351 && y == 7'd235) || (x == 7'd634 && y == 7'd57) ||
		(x == 7'd343 && y == 179) || (x == 7'd582 && y == 628) || (x == 7'd404 && y == 7'd260) ||
		(x == 7'd270 && y == 577) || (x == 562 && y == 199) || (x == 7'd144 && y == 451) ||
		(x == 330 && y == 7'd123) || (x == 7'd111 && y == 94) || (x == 7'd532 && y == 110) ||
		(x == 244 && y == 7'd19) || (x == 7'd64 && y == 71) || (x == 7'd154 && y == 7'd483) ||
		(x == 7'd111 && y == 161) || (x == 7'd489 && y == 204) || (x == 7'd389 && y == 73) ||
		(x == 357 && y == 7'd346) || (x == 579 && y == 263) || (x == 70 && y == 7'd564) ||
		(x == 7'd461 && y == 81) || (x == 7'd534 && y == 7'd80) || (x == 366 && y == 616) ||
		(x == 7'd438 && y == 7'd637) || (x == 7'd9 && y == 526) || (x == 547 && y == 7'd523) ||
		(x == 369 && y == 292) || (x == 7'd226 && y == 7'd489) || (x == 210 && y == 469) ||
		(x == 137 && y == 175) || (x == 435 && y == 245) || (x == 7'd442 && y == 7'd622) ||
		(x == 7'd79 && y == 7'd598) || (x == 495 && y == 7'd258) || (x == 7'd276 && y == 7'd283) ||
		(x == 7'd315 && y == 301) || (x == 7'd7 && y == 609) || (x == 144 && y == 7'd190) ||
		(x == 225 && y == 368) || (x == 7'd476 && y == 7'd240) || (x == 505 && y == 441) ||
		(x == 7'd323 && y == 7'd210) || (x == 545 && y == 7'd300) || (x == 7'd267 && y == 7'd442) ||
		(x == 7'd370 && y == 495) || (x == 492 && y == 482) || (x == 7'd427 && y == 7'd523) ||
		(x == 373 && y == 618) || (x == 7'd189 && y == 122) || (x == 7'd455 && y == 7'd306) ||
		(x == 7'd353 && y == 7'd144) || (x == 7'd299 && y == 7'd392) || (x == 7'd609 && y == 7'd439) ||
		(x == 551 && y == 7'd17) || (x == 7'd209 && y == 548) || (x == 19 && y == 7'd620) ||
		(x == 7'd160 && y == 7'd300) || (x == 7'd116 && y == 148) || (x == 7'd480 && y == 7'd238) ||
		(x == 108 && y == 7'd147) || (x == 7'd288 && y == 519) || (x == 296 && y == 7'd149) ||
		(x == 7'd169 && y == 7'd223) || (x == 7'd373 && y == 534) || (x == 241 && y == 417) ||
		(x == 348 && y == 472) || (x == 7'd342 && y == 285) || (x == 335 && y == 7'd625) ||
		(x == 175 && y == 367) || (x == 449 && y == 7'd351) || (x == 7'd287 && y == 7'd402) ||
		(x == 7'd614 && y == 7'd275) || (x == 486 && y == 426) || (x == 636 && y == 636) ||
		(x == 7'd132 && y == 7'd452) || (x == 7'd319 && y == 7'd134) || (x == 607 && y == 7'd183) ||
		(x == 7'd268 && y == 7'd502) || (x == 550 && y == 436) || (x == 7'd320 && y == 7'd551) ||
		(x == 195 && y == 7'd540) || (x == 7'd132 && y == 7'd306) || (x == 7'd186 && y == 7'd580) ||
		(x == 7'd275 && y == 7'd155) || (x == 7'd272 && y == 319) || (x == 7'd623 && y == 7'd310) ||
		(x == 7'd250 && y == 7'd634) || (x == 280 && y == 7'd454) || (x == 310 && y == 7'd557) ||
		(x == 556 && y == 131) || (x == 298 && y == 7'd411) || (x == 7'd264 && y == 231) ||
		(x == 7'd158 && y == 7'd413) || (x == 7'd363 && y == 28) || (x == 344 && y == 318) ||
		(x == 7'd574 && y == 582) || (x == 7'd140 && y == 181) || (x == 7'd579 && y == 7'd593) ||
		(x == 131 && y == 7'd111) || (x == 7'd80 && y == 325) || (x == 7'd444 && y == 7'd475) ||
		(x == 7'd253 && y == 7'd429) || (x == 306 && y == 7'd550) || (x == 178 && y == 7'd539) ||
		(x == 526 && y == 504) || (x == 7'd503 && y == 455) || (x == 7'd530 && y == 55) ||
		(x == 7'd523 && y == 87) || (x == 466 && y == 7'd262) || (x == 526 && y == 141) ||
		(x == 7'd211 && y == 7'd388) || (x == 7'd479 && y == 7'd213) || (x == 7'd118 && y == 369) ||
		(x == 7'd80 && y == 364) || (x == 585 && y == 245) || (x == 558 && y == 7'd246) ||
		(x == 7'd519 && y == 7'd259) || (x == 7'd336 && y == 7'd366) || (x == 7'd383 && y == 65) ||
		(x == 598 && y == 7'd439) || (x == 207 && y == 627) || (x == 298 && y == 7'd532) ||
		(x == 379 && y == 7'd421) || (x == 7'd244 && y == 14) || (x == 7'd263 && y == 7'd181) ||
		(x == 7'd569 && y == 7'd401) || (x == 147 && y == 7'd210) || (x == 20 && y == 7'd415) ||
		(x == 472 && y == 7'd145) || (x == 241 && y == 7'd246) || (x == 7'd618 && y == 534) ||
		(x == 7'd430 && y == 7'd140) || (x == 7'd297 && y == 7'd599) || (x == 631 && y == 153) ||
		(x == 7'd479 && y == 7'd336) || (x == 348 && y == 7'd30) || (x == 7'd625 && y == 7'd310) ||
		(x == 7'd186 && y == 7'd346) || (x == 7'd518 && y == 7'd353) || (x == 7'd267 && y == 7'd527) ||
		(x == 474 && y == 7'd567) || (x == 7'd244 && y == 7'd457) || (x == 7'd534 && y == 7'd139) ||
		(x == 7'd388 && y == 7'd581) || (x == 7'd355 && y == 7'd272) || (x == 7'd369 && y == 7'd239) ||
		(x == 478 && y == 7'd542) || (x == 13 && y == 7'd298) || (x == 7'd335 && y == 7'd20) ||
		(x == 470 && y == 7'd158) || (x == 7'd268 && y == 528) || (x == 7'd296 && y == 406) ||
		(x == 7'd418 && y == 7'd470) || (x == 381 && y == 170) || (x == 485 && y == 7'd86) ||
		(x == 7'd399 && y == 7'd172) || (x == 432 && y == 7'd20) || (x == 7'd242 && y == 7'd94) ||
		(x == 7'd117 && y == 7'd600) || (x == 7'd382 && y == 257) || (x == 494 && y == 596) ||
		(x == 7'd441 && y == 7'd399) || (x == 7'd551 && y == 7'd629) || (x == 542 && y == 609) ||
		(x == 374 && y == 7'd24) || (x == 536 && y == 7'd220) || (x == 7'd338 && y == 586) ||
		(x == 130 && y == 421) || (x == 366 && y == 7'd468) || (x == 220 && y == 216) ||
		(x == 7'd41 && y == 98) || (x == 7'd165 && y == 7'd245) || (x == 7'd576 && y == 7'd249) ||
		(x == 7'd433 && y == 7'd399) || (x == 185 && y == 230) || (x == 6 && y == 7'd238) ||
		(x == 7'd302 && y == 7'd635) || (x == 7'd437 && y == 7'd253) || (x == 611 && y == 174) ||
		(x == 278 && y == 7'd210) || (x == 7'd488 && y == 638) || (x == 89 && y == 7'd380) ||
		(x == 218 && y == 535) || (x == 131 && y == 7'd60) || (x == 479 && y == 7'd305) ||
		(x == 7'd162 && y == 7'd228) || (x == 367 && y == 131) || (x == 7'd269 && y == 7'd148) ||
		(x == 7'd450 && y == 96) || (x == 87 && y == 7'd589) || (x == 7'd44 && y == 7'd326) ||
		(x == 7'd612 && y == 7'd424) || (x == 503 && y == 7'd331) || (x == 7'd548 && y == 7'd157) ||
		(x == 403 && y == 7'd369) || (x == 397 && y == 130) || (x == 435 && y == 167) ||
		(x == 331 && y == 7'd235) || (x == 7'd448 && y == 483) || (x == 7'd126 && y == 233) ||
		(x == 142 && y == 345) || (x == 7'd630 && y == 7'd478) || (x == 7'd407 && y == 7'd410) ||
		(x == 348 && y == 7'd241) || (x == 356 && y == 7'd227) || (x == 7'd352 && y == 17) ||
		(x == 7'd507 && y == 7'd274) || (x == 7'd187 && y == 183) || (x == 7'd370 && y == 7'd448) ||
		(x == 143 && y == 486) || (x == 7'd592 && y == 7'd121) || (x == 561 && y == 7'd231) ||
		(x == 7'd522 && y == 7'd385) || (x == 7'd363 && y == 7'd429) || (x == 7'd105 && y == 7'd276) ||
		(x == 7'd599 && y == 7'd402) || (x == 537 && y == 7'd382) || (x == 456 && y == 347) ||
		(x == 276 && y == 313) || (x == 63 && y == 7'd199) || (x == 7'd171 && y == 487) ||
		(x == 581 && y == 505) || (x == 577 && y == 634) || (x == 7'd145 && y == 7'd369) ||
		(x == 626 && y == 7'd605) || (x == 7'd339 && y == 7'd209) || (x == 335 && y == 7'd555) ||
		(x == 250 && y == 7'd406) || (x == 7'd27 && y == 542) || (x == 7'd503 && y == 63) ||
		(x == 7 && y == 7'd591) || (x == 7'd578 && y == 7'd107) || (x == 7'd621 && y == 7'd27) ||
		(x == 549 && y == 7'd151) || (x == 7'd632 && y == 260) || (x == 7'd543 && y == 638) ||
		(x == 7'd413 && y == 455) || (x == 562 && y == 7'd46) || (x == 7'd465 && y == 7'd380) ||
		(x == 192 && y == 7'd578) || (x == 154 && y == 173) || (x == 7'd71 && y == 7'd542) ||
		(x == 7'd380 && y == 188) || (x == 7'd620 && y == 470) || (x == 7'd215 && y == 513) ||
		(x == 47 && y == 7'd190) || (x == 7'd475 && y == 525) || (x == 242 && y == 314) ||
		(x == 7'd450 && y == 612) || (x == 40 && y == 7'd264) || (x == 267 && y == 505) ||
		(x == 7'd351 && y == 7'd525) || (x == 603 && y == 7'd78) || (x == 21 && y == 7'd462) ||
		(x == 196 && y == 7'd204) || (x == 558 && y == 7'd287) || (x == 7'd362 && y == 7'd635) ||
		(x == 491 && y == 528) || (x == 7'd339 && y == 7'd245) || (x == 7'd563 && y == 157) ||
		(x == 7'd65 && y == 214) || (x == 145 && y == 7'd380) || (x == 7'd427 && y == 224) ||
		(x == 227 && y == 7'd439) || (x == 7'd590 && y == 44) || (x == 7'd625 && y == 7'd582) ||
		(x == 7'd601 && y == 7'd370) || (x == 7'd177 && y == 7'd526) || (x == 452 && y == 596) ||
		(x == 127 && y == 7'd175) || (x == 186 && y == 223) || (x == 224 && y == 7'd539) ||
		(x == 178 && y == 7'd478) || (x == 7'd455 && y == 608) || (x == 7'd573 && y == 7'd259) ||
		(x == 7'd436 && y == 7'd527) || (x == 7'd57 && y == 384) || (x == 7'd462 && y == 543) ||
		(x == 447 && y == 544) || (x == 7'd141 && y == 235) || (x == 504 && y == 541) ||
		(x == 7'd112 && y == 7'd377) || (x == 7'd378 && y == 7'd505) || (x == 7'd511 && y == 7'd228) ||
		(x == 302 && y == 399) || (x == 7'd254 && y == 7'd325) || (x == 7'd100 && y == 7'd149) ||
		(x == 450 && y == 219) || (x == 7'd366 && y == 7'd401) || (x == 7'd231 && y == 7'd638) ||
		(x == 7'd251 && y == 7'd143) || (x == 342 && y == 7'd366) || (x == 426 && y == 7'd47) ||
		(x == 7'd421 && y == 202) || (x == 7'd63 && y == 308) || (x == 7'd21 && y == 340) ||
		(x == 402 && y == 375) || (x == 7'd245 && y == 7'd583) || (x == 485 && y == 7'd493) ||
		(x == 7'd556 && y == 506) || (x == 7'd136 && y == 7'd75) || (x == 7'd282 && y == 606) ||
		(x == 7'd223 && y == 126) || (x == 7'd563 && y == 7'd403) || (x == 7'd498 && y == 327) ||
		(x == 7'd527 && y == 112) || (x == 301 && y == 280) || (x == 7'd181 && y == 525) ||
		(x == 627 && y == 544) || (x == 7'd223 && y == 7'd46) || (x == 7'd394 && y == 213) ||
		(x == 7'd379 && y == 573) || (x == 72 && y == 7'd133) || (x == 417 && y == 217) ||
		(x == 601 && y == 7'd480) || (x == 7'd164 && y == 7'd627) || (x == 7'd289 && y == 62) ||
		(x == 296 && y == 592) || (x == 448 && y == 321) || (x == 278 && y == 627) ||
		(x == 7'd468 && y == 481) || (x == 477 && y == 287) || (x == 7'd216 && y == 7'd262) ||
		(x == 7'd352 && y == 565) || (x == 7'd290 && y == 7'd247) || (x == 227 && y == 7'd58) ||
		(x == 7'd46 && y == 7'd552) || (x == 491 && y == 411) || (x == 431 && y == 343) ||
		(x == 366 && y == 365) || (x == 7'd260 && y == 7'd364) || (x == 7'd504 && y == 7'd459) ||
		(x == 7'd442 && y == 7'd377) || (x == 7'd495 && y == 7'd158) || (x == 508 && y == 205) ||
		(x == 270 && y == 7'd553) || (x == 478 && y == 7'd542) || (x == 7'd282 && y == 7'd201) ||
		(x == 7'd447 && y == 7'd558) || (x == 7'd166 && y == 7'd198) || (x == 139 && y == 485) ||
		(x == 590 && y == 7'd320) || (x == 528 && y == 359) || (x == 7'd565 && y == 591) ||
		(x == 446 && y == 543) || (x == 7'd223 && y == 277) || (x == 7'd60 && y == 153) ||
		(x == 7'd112 && y == 7'd423) || (x == 7'd490 && y == 7'd555) || (x == 7'd589 && y == 7'd426) ||
		(x == 343 && y == 7'd154) || (x == 177 && y == 191) || (x == 7'd135 && y == 7'd385) ||
		(x == 7'd178 && y == 7'd254) || (x == 7'd65 && y == 7'd570) || (x == 7'd473 && y == 7'd10) ||
		(x == 414 && y == 7'd28) || (x == 576 && y == 7'd577) || (x == 7'd262 && y == 265) ||
		(x == 387 && y == 453) || (x == 7'd288 && y == 255) || (x == 267 && y == 152) ||
		(x == 7'd386 && y == 7'd519) || (x == 549 && y == 7'd624) || (x == 7'd626 && y == 7'd141) ||
		(x == 7'd364 && y == 569) || (x == 7'd639 && y == 7'd26) || (x == 7'd112 && y == 553) ||
		(x == 383 && y == 7'd453) || (x == 7'd530 && y == 7'd340) || (x == 141 && y == 7'd555) ||
		(x == 7'd102 && y == 7'd182) || (x == 602 && y == 527) || (x == 7'd614 && y == 7'd466) ||
		(x == 369 && y == 168) || (x == 7'd523 && y == 7'd575) || (x == 303 && y == 178) ||
		(x == 7'd130 && y == 7'd264) || (x == 620 && y == 7'd198) || (x == 540 && y == 144) ||
		(x == 443 && y == 7'd428) || (x == 545 && y == 534) || (x == 273 && y == 7'd311) ||
		(x == 7'd128 && y == 539) || (x == 593 && y == 202) || (x == 7'd445 && y == 405) ||
		(x == 7'd345 && y == 7'd583) || (x == 180 && y == 7'd304) || (x == 7'd576 && y == 7'd169) ||
		(x == 7'd428 && y == 7'd460) || (x == 7'd570 && y == 202) || (x == 7'd35 && y == 414) ||
		(x == 437 && y == 7'd119) || (x == 7'd61 && y == 606) || (x == 7'd557 && y == 611) ||
		(x == 616 && y == 226) || (x == 7'd291 && y == 7'd204) || (x == 304 && y == 7'd358) ||
		(x == 7'd160 && y == 7'd85) || (x == 7'd16 && y == 7'd534) || (x == 7'd221 && y == 7'd174) ||
		(x == 7'd582 && y == 498) || (x == 481 && y == 616) || (x == 7'd555 && y == 81) ||
		(x == 163 && y == 7'd401) || (x == 178 && y == 369) || (x == 187 && y == 7'd338) ||
		(x == 7'd319 && y == 455) || (x == 371 && y == 7'd192) || (x == 7'd44 && y == 266) ||
		(x == 7'd555 && y == 503) || (x == 308 && y == 450) || (x == 7'd616 && y == 7'd623) ||
		(x == 433 && y == 7'd617) || (x == 7'd423 && y == 7'd486) || (x == 7'd439 && y == 7'd466) ||
		(x == 75 && y == 7'd146) || (x == 7'd371 && y == 7'd521) || (x == 7'd623 && y == 7'd629) ||
		(x == 7'd410 && y == 7'd225) || (x == 7'd622 && y == 7'd178) || (x == 170 && y == 366) ||
		(x == 334 && y == 638) || (x == 129 && y == 7'd395) || (x == 195 && y == 617) ||
		(x == 7'd516 && y == 7'd564) || (x == 526 && y == 254) || (x == 301 && y == 151) ||
		(x == 544 && y == 504) || (x == 559 && y == 7'd343) || (x == 7'd358 && y == 7'd623) ||
		(x == 7'd632 && y == 7'd235) || (x == 7'd358 && y == 7'd404) || (x == 7'd196 && y == 7'd39) ||
		(x == 441 && y == 536) || (x == 7'd274 && y == 7'd111) || (x == 7'd211 && y == 7'd179) ||
		(x == 7'd582 && y == 7'd400) || (x == 366 && y == 526) || (x == 304 && y == 7'd119) ||
		(x == 82 && y == 7'd243) || (x == 349 && y == 433) || (x == 7'd193 && y == 7'd354) ||
		(x == 239 && y == 483) || (x == 251 && y == 446) || (x == 254 && y == 596) ||
		(x == 7'd334 && y == 188) || (x == 180 && y == 565) || (x == 7'd574 && y == 446) ||
		(x == 231 && y == 7'd315) || (x == 7'd201 && y == 7'd610) || (x == 7'd621 && y == 639) ||
		(x == 635 && y == 327) || (x == 7'd368 && y == 7'd241) || (x == 7'd213 && y == 495) ||
		(x == 7'd161 && y == 7'd512) || (x == 506 && y == 560) || (x == 7'd41 && y == 9) ||
		(x == 7'd511 && y == 7'd281) || (x == 7'd568 && y == 7'd71) || (x == 7'd47 && y == 7'd11) ||
		(x == 149 && y == 7'd395) || (x == 566 && y == 7'd159) || (x == 142 && y == 7'd77) ||
		(x == 608 && y == 131) || (x == 7'd557 && y == 7'd264) || (x == 7'd270 && y == 7'd58) ||
		(x == 7'd392 && y == 7'd420) || (x == 325 && y == 257) || (x == 7'd550 && y == 7'd628) ||
		(x == 249 && y == 7'd569) || (x == 7'd541 && y == 583) || (x == 7'd426 && y == 7'd132) ||
		(x == 455 && y == 7'd162) || (x == 7'd200 && y == 582) || (x == 583 && y == 379) ||
		(x == 7'd225 && y == 7'd270) || (x == 7'd494 && y == 7'd347) || (x == 434 && y == 7'd87) ||
		(x == 7'd144 && y == 35) || (x == 7'd497 && y == 7'd583) || (x == 59 && y == 7'd627) ||
		(x == 259 && y == 256) || (x == 7'd382 && y == 7'd502) || (x == 246 && y == 547) ||
		(x == 467 && y == 608) || (x == 567 && y == 7'd533) || (x == 61 && y == 7'd141) ||
		(x == 233 && y == 287) || (x == 121 && y == 7'd164) || (x == 592 && y == 538) ||
		(x == 7'd214 && y == 7'd550) || (x == 145 && y == 7'd224) || (x == 7'd298 && y == 259) ||
		(x == 380 && y == 424) || (x == 139 && y == 562) || (x == 271 && y == 232) ||
		(x == 451 && y == 399) || (x == 168 && y == 144) || (x == 7'd540 && y == 7'd269) ||
		(x == 7'd577 && y == 7'd137) || (x == 240 && y == 7'd247) || (x == 7'd199 && y == 7'd625) ||
		(x == 7'd62 && y == 620) || (x == 508 && y == 590) || (x == 7'd193 && y == 7'd86) ||
		(x == 7'd265 && y == 7'd461) || (x == 7'd573 && y == 7'd134) || (x == 7'd598 && y == 7'd503) ||
		(x == 7'd478 && y == 262) || (x == 50 && y == 14) || (x == 377 && y == 191) ||
		(x == 7'd61 && y == 41) || (x == 265 && y == 7'd53) || (x == 336 && y == 144) ||
		(x == 621 && y == 7'd288) || (x == 620 && y == 261) || (x == 7'd352 && y == 387) ||
		(x == 7'd130 && y == 522) || (x == 7'd344 && y == 7'd347) || (x == 131 && y == 161) ||
		(x == 7'd439 && y == 192) || (x == 7'd373 && y == 196) || (x == 7'd632 && y == 7'd393) ||
		(x == 414 && y == 7'd120) || (x == 7'd536 && y == 255) || (x == 318 && y == 565) ||
		(x == 7'd41 && y == 565) || (x == 179 && y == 530) || (x == 7'd498 && y == 7'd393) ||
		(x == 605 && y == 294) || (x == 7'd462 && y == 7'd276) || (x == 7'd619 && y == 7'd47) ||
		(x == 7'd580 && y == 7'd202) || (x == 515 && y == 577) || (x == 7'd217 && y == 7'd132) ||
		(x == 501 && y == 427) || (x == 19 && y == 7'd518) || (x == 7'd533 && y == 7'd178) ||
		(x == 383 && y == 7'd73) || (x == 342 && y == 239) || (x == 560 && y == 7'd24) ||
		(x == 7'd242 && y == 636) || (x == 331 && y == 303) || (x == 340 && y == 313) ||
		(x == 7'd425 && y == 73) || (x == 227 && y == 476) || (x == 7'd409 && y == 7'd560) ||
		(x == 7'd398 && y == 569) || (x == 7'd191 && y == 319) || (x == 273 && y == 394) ||
		(x == 7'd158 && y == 7'd586) || (x == 409 && y == 7'd528) || (x == 254 && y == 7'd454) ||
		(x == 7'd428 && y == 7'd594) || (x == 7'd465 && y == 321) || (x == 555 && y == 596) ||
		(x == 274 && y == 7'd196) || (x == 7'd538 && y == 7'd437) || (x == 7'd58 && y == 280) ||
		(x == 7'd438 && y == 189) || (x == 215 && y == 7'd116) || (x == 7'd545 && y == 435) ||
		(x == 181 && y == 7'd480) || (x == 7'd426 && y == 324) || (x == 7'd398 && y == 575) ||
		(x == 7'd177 && y == 7'd363) || (x == 527 && y == 352) || (x == 417 && y == 7'd344) ||
		(x == 7'd266 && y == 7'd23) || (x == 504 && y == 539) || (x == 359 && y == 7'd414) ||
		(x == 7'd634 && y == 7'd211) || (x == 617 && y == 335) || (x == 450 && y == 429) ||
		(x == 597 && y == 506) || (x == 7'd20 && y == 7'd206) || (x == 308 && y == 244) ||
		(x == 7'd486 && y == 7'd561) || (x == 498 && y == 170) || (x == 576 && y == 385) ||
		(x == 7'd615 && y == 1) || (x == 7'd277 && y == 7'd268) || (x == 58 && y == 7'd628) ||
		(x == 7'd381 && y == 7'd143) || (x == 7'd62 && y == 367) || (x == 515 && y == 571) ||
		(x == 454 && y == 7'd560) || (x == 303 && y == 7'd476) || (x == 7'd549 && y == 7'd289) ||
		(x == 174 && y == 7'd183) || (x == 118 && y == 7'd8) || (x == 7'd316 && y == 7'd600) ||
		(x == 332 && y == 7'd92) || (x == 578 && y == 196) || (x == 7'd596 && y == 385) ||
		(x == 7'd162 && y == 7'd64) || (x == 7'd446 && y == 7'd101) || (x == 613 && y == 7'd27) ||
		(x == 180 && y == 7'd332) || (x == 7'd22 && y == 489) || (x == 7'd448 && y == 347) ||
		(x == 386 && y == 7'd490) || (x == 7'd134 && y == 7'd635) || (x == 137 && y == 7'd367) ||
		(x == 322 && y == 296) || (x == 7'd592 && y == 162) || (x == 307 && y == 7'd252) ||
		(x == 492 && y == 418) || (x == 7'd316 && y == 250) || (x == 7'd78 && y == 403) ||
		(x == 7'd258 && y == 586) || (x == 388 && y == 292) || (x == 7'd445 && y == 7'd246) ||
		(x == 7'd209 && y == 7'd29) || (x == 7'd297 && y == 346) || (x == 14 && y == 7'd450) ||
		(x == 7'd470 && y == 536) || (x == 7'd84 && y == 248) || (x == 7'd111 && y == 7'd171) ||
		(x == 7'd266 && y == 7'd547) || (x == 604 && y == 7'd247) || (x == 7'd599 && y == 7'd136) ||
		(x == 234 && y == 375) || (x == 7'd111 && y == 7'd324) || (x == 352 && y == 523) ||
		(x == 7'd468 && y == 7'd284) || (x == 7'd410 && y == 7'd301) || (x == 7'd347 && y == 7'd482) ||
		(x == 277 && y == 7'd596) || (x == 7'd581 && y == 13) || (x == 7'd271 && y == 7'd189) ||
		(x == 566 && y == 436) || (x == 256 && y == 7'd491) || (x == 7'd366 && y == 273) ||
		(x == 7'd519 && y == 7'd590) || (x == 7'd137 && y == 7'd403) || (x == 488 && y == 7'd357) ||
		(x == 7'd605 && y == 554) || (x == 7'd168 && y == 7'd491) || (x == 7'd92 && y == 7'd239) ||
		(x == 7'd627 && y == 217) || (x == 7'd161 && y == 627) || (x == 450 && y == 637) ||
		(x == 7'd231 && y == 7'd626) || (x == 361 && y == 7'd412) || (x == 508 && y == 7'd500) ||
		(x == 398 && y == 320) || (x == 7'd575 && y == 7'd166) || (x == 7'd476 && y == 7'd177) ||
		(x == 120 && y == 7'd379) || (x == 191 && y == 513) || (x == 7'd620 && y == 328) ||
		(x == 147 && y == 606) || (x == 7'd103 && y == 7'd378) || (x == 580 && y == 7'd461) ||
		(x == 240 && y == 7'd29) || (x == 376 && y == 7'd0) || (x == 7'd285 && y == 511) ||
		(x == 7'd545 && y == 145) || (x == 7'd192 && y == 7'd340) || (x == 7'd269 && y == 601) ||
		(x == 409 && y == 494) || (x == 7'd393 && y == 7'd631) || (x == 7'd368 && y == 322) ||
		(x == 312 && y == 253) || (x == 7'd237 && y == 7'd220) || (x == 62 && y == 7'd295) ||
		(x == 7'd255 && y == 7'd435) || (x == 7'd507 && y == 245) || (x == 7'd149 && y == 603) ||
		(x == 7'd316 && y == 84) || (x == 385 && y == 588) || (x == 7'd614 && y == 7'd48) ||
		(x == 7'd283 && y == 7'd556) || (x == 221 && y == 381) || (x == 470 && y == 7'd45) ||
		(x == 166 && y == 7'd562) || (x == 7'd228 && y == 429) || (x == 229 && y == 7'd88) ||
		(x == 7'd254 && y == 248) || (x == 473 && y == 357) || (x == 510 && y == 7'd239) ||
		(x == 534 && y == 7'd332) || (x == 374 && y == 350) || (x == 7'd575 && y == 213) ||
		(x == 373 && y == 247) || (x == 7'd163 && y == 7'd574) || (x == 7'd262 && y == 7'd196) ||
		(x == 7'd378 && y == 7'd619) || (x == 7'd315 && y == 605) || (x == 596 && y == 7'd386) ||
		(x == 7'd612 && y == 7'd176) || (x == 7'd520 && y == 7'd58) || (x == 125 && y == 7'd229) ||
		(x == 7'd61 && y == 162) || (x == 7'd33 && y == 7'd247) || (x == 621 && y == 7'd386) ||
		(x == 223 && y == 388) || (x == 7'd534 && y == 7'd582) || (x == 289 && y == 183) ||
		(x == 7'd593 && y == 7'd251) || (x == 419 && y == 7'd161) || (x == 7'd534 && y == 632) ||
		(x == 7'd594 && y == 258) || (x == 7'd400 && y == 7'd531) || (x == 7'd149 && y == 7'd325) ||
		(x == 413 && y == 7'd13) || (x == 7'd19 && y == 7'd280) || (x == 7'd416 && y == 7'd423) ||
		(x == 7'd405 && y == 7'd252) || (x == 7'd430 && y == 346) || (x == 7'd167 && y == 7'd526) ||
		(x == 7'd325 && y == 7'd329) || (x == 7'd209 && y == 269) || (x == 495 && y == 433) ||
		(x == 7'd633 && y == 7'd540) || (x == 7'd0 && y == 299) || (x == 139 && y == 7'd563) ||
		(x == 7'd155 && y == 7'd350) || (x == 565 && y == 7'd226) || (x == 549 && y == 7'd612) ||
		(x == 7'd305 && y == 7'd514) || (x == 7'd6 && y == 247) || (x == 7'd391 && y == 7'd560) ||
		(x == 7'd9 && y == 213) || (x == 291 && y == 7'd342) || (x == 424 && y == 298) ||
		(x == 293 && y == 7'd333) || (x == 7'd415 && y == 7'd286) || (x == 7'd362 && y == 596) ||
		(x == 7'd313 && y == 7'd377) || (x == 7'd414 && y == 68) || (x == 522 && y == 7'd298) ||
		(x == 7'd391 && y == 7'd289) || (x == 7'd532 && y == 261) || (x == 7'd635 && y == 7'd414) ||
		(x == 7'd349 && y == 533) || (x == 7'd239 && y == 281) || (x == 384 && y == 7'd43) ||
		(x == 131 && y == 492) || (x == 7'd465 && y == 418) || (x == 57 && y == 7'd254) ||
		(x == 7'd392 && y == 7'd299) || (x == 303 && y == 250) || (x == 244 && y == 551) ||
		(x == 7'd496 && y == 7'd630) || (x == 7'd76 && y == 303) || (x == 7'd322 && y == 291) ||
		(x == 468 && y == 7'd521) || (x == 279 && y == 7'd13) || (x == 7'd442 && y == 7'd143) ||
		(x == 7'd491 && y == 7'd373) || (x == 7'd588 && y == 50) || (x == 189 && y == 7'd186) ||
		(x == 7'd224 && y == 7'd293) || (x == 7'd425 && y == 7'd432) || (x == 33 && y == 7'd346) ||
		(x == 7'd16 && y == 7'd24) || (x == 7'd38 && y == 7'd384) || (x == 151 && y == 321) ||
		(x == 7'd242 && y == 7'd70) || (x == 246 && y == 366) || (x == 200 && y == 7'd157) ||
		(x == 7'd26 && y == 7'd545) || (x == 600 && y == 7'd275) || (x == 7'd130 && y == 7'd232) ||
		(x == 329 && y == 7'd430) || (x == 7'd586 && y == 514) || (x == 7'd409 && y == 572) ||
		(x == 71 && y == 7'd525) || (x == 121 && y == 7'd554) || (x == 474 && y == 435) ||
		(x == 178 && y == 342) || (x == 7'd126 && y == 7'd375) || (x == 296 && y == 7'd201) ||
		(x == 7'd154 && y == 7'd460) || (x == 7'd422 && y == 7'd4) || (x == 7'd16 && y == 525) ||
		(x == 213 && y == 7'd237) || (x == 521 && y == 420) || (x == 7'd67 && y == 7'd177) ||
		(x == 7'd285 && y == 7'd465) || (x == 7'd458 && y == 566) || (x == 7'd228 && y == 7'd300) ||
		(x == 7'd444 && y == 7'd272) || (x == 7'd130 && y == 7'd540) || (x == 7'd450 && y == 7'd432) ||
		(x == 210 && y == 528) || (x == 159 && y == 7'd169) || (x == 197 && y == 7'd359) ||
		(x == 283 && y == 7'd146) || (x == 468 && y == 7'd566) || (x == 7'd378 && y == 7'd554) ||
		(x == 7'd634 && y == 7'd487) || (x == 7'd283 && y == 214) || (x == 7'd116 && y == 7'd624) ||
		(x == 7'd363 && y == 7'd512) || (x == 7'd633 && y == 7'd39) || (x == 147 && y == 7'd436) ||
		(x == 7'd459 && y == 7'd172) || (x == 264 && y == 7'd566) || (x == 431 && y == 7'd306) ||
		(x == 7'd420 && y == 7'd483) || (x == 486 && y == 606) || (x == 7'd612 && y == 126) ||
		(x == 7'd612 && y == 7'd308) || (x == 8 && y == 7'd605) || (x == 220 && y == 7'd365) ||
		(x == 7'd4 && y == 7'd352) || (x == 359 && y == 7'd250) || (x == 7'd583 && y == 7'd207) ||
		(x == 453 && y == 7'd260) || (x == 7'd242 && y == 369) || (x == 7'd474 && y == 7'd134) ||
		(x == 7'd5 && y == 7'd538) || (x == 7'd99 && y == 7'd621) || (x == 7'd442 && y == 7'd581) ||
		(x == 254 && y == 143) || (x == 7'd532 && y == 7'd43) || (x == 7'd282 && y == 565) ||
		(x == 292 && y == 7'd9) || (x == 578 && y == 282) || (x == 386 && y == 7'd307) ||
		(x == 474 && y == 574) || (x == 583 && y == 7'd210) || (x == 7'd246 && y == 7'd467) ||
		(x == 114 && y == 7'd479) || (x == 7'd609 && y == 597) || (x == 7'd200 && y == 334) ||
		(x == 7'd476 && y == 7'd243) || (x == 7'd306 && y == 183) || (x == 7'd575 && y == 550) ||
		(x == 7'd495 && y == 7'd539) || (x == 177 && y == 159) || (x == 7'd633 && y == 7'd159) ||
		(x == 152 && y == 401) || (x == 7'd453 && y == 618) || (x == 480 && y == 7'd120) ||
		(x == 219 && y == 7'd319) || (x == 7'd260 && y == 7'd477) || (x == 7'd397 && y == 7'd468) ||
		(x == 28 && y == 7'd526) || (x == 375 && y == 7'd182) || (x == 7'd516 && y == 7'd141) ||
		(x == 297 && y == 381) || (x == 496 && y == 326) || (x == 7'd159 && y == 7'd15) ||
		(x == 7'd412 && y == 7'd516) || (x == 7'd241 && y == 7'd478) || (x == 355 && y == 423) ||
		(x == 7'd463 && y == 7'd230) || (x == 7'd571 && y == 15) || (x == 7'd95 && y == 329) ||
		(x == 7'd370 && y == 7'd456) || (x == 131 && y == 7'd419) || (x == 7'd63 && y == 448) ||
		(x == 184 && y == 435) || (x == 7'd446 && y == 332) || (x == 236 && y == 7'd92) ||
		(x == 7'd530 && y == 277) || (x == 273 && y == 7'd268) || (x == 7'd474 && y == 7'd561) ||
		(x == 286 && y == 7'd441) || (x == 7'd331 && y == 537) || (x == 215 && y == 7'd24) ||
		(x == 7'd450 && y == 7'd379) || (x == 7'd542 && y == 7'd119) || (x == 7'd382 && y == 7'd436) ||
		(x == 7'd434 && y == 7'd459) || (x == 590 && y == 7'd155) || (x == 7'd505 && y == 7'd399) ||
		(x == 519 && y == 7'd316) || (x == 242 && y == 7'd88) || (x == 7'd18 && y == 7'd209) ||
		(x == 388 && y == 366) || (x == 7'd623 && y == 118) || (x == 7'd402 && y == 7'd389) ||
		(x == 505 && y == 151) || (x == 261 && y == 7'd546) || (x == 7'd533 && y == 7'd133) ||
		(x == 7'd417 && y == 359) || (x == 7'd308 && y == 7'd403) || (x == 7'd374 && y == 7'd447) ||
		(x == 576 && y == 393) || (x == 300 && y == 622) || (x == 605 && y == 7'd65) ||
		(x == 7'd508 && y == 7'd537) || (x == 7'd103 && y == 204) || (x == 607 && y == 7'd402) ||
		(x == 329 && y == 7'd142) || (x == 483 && y == 235) || (x == 577 && y == 7'd70) ||
		(x == 251 && y == 294) || (x == 7'd229 && y == 7'd240) || (x == 228 && y == 522) ||
		(x == 7'd99 && y == 283) || (x == 586 && y == 7'd582) || (x == 7'd33 && y == 617) ||
		(x == 476 && y == 7'd531) || (x == 545 && y == 503) || (x == 512 && y == 7'd270) ||
		(x == 7'd362 && y == 134) || (x == 7'd184 && y == 7'd513) || (x == 7'd379 && y == 7'd362) ||
		(x == 158 && y == 7'd627) || (x == 361 && y == 7'd448) || (x == 7'd214 && y == 7'd79) ||
		(x == 19 && y == 7'd197) || (x == 7'd126 && y == 419) || (x == 79 && y == 7'd251) ||
		(x == 495 && y == 489) || (x == 7'd48 && y == 395) || (x == 7'd468 && y == 7'd389) ||
		(x == 599 && y == 7'd476) || (x == 7'd33 && y == 7'd529) || (x == 7'd529 && y == 7'd410) ||
		(x == 213 && y == 7'd80) || (x == 7'd376 && y == 7'd361) || (x == 7'd147 && y == 170) ||
		(x == 246 && y == 224) || (x == 414 && y == 601) || (x == 7'd255 && y == 7'd500) ||
		(x == 7'd413 && y == 7'd256) || (x == 7'd81 && y == 491) || (x == 7'd138 && y == 7'd315) ||
		(x == 7'd142 && y == 7'd497) || (x == 7'd503 && y == 7'd78) || (x == 404 && y == 207) ||
		(x == 7'd373 && y == 7'd492) || (x == 7'd613 && y == 7'd262) || (x == 7'd308 && y == 516) ||
		(x == 7'd324 && y == 75) || (x == 473 && y == 7'd623) || (x == 123 && y == 7'd122) ||
		(x == 7'd342 && y == 7'd371) || (x == 113 && y == 7'd260) || (x == 7'd369 && y == 7'd144) ||
		(x == 556 && y == 548) || (x == 432 && y == 566) || (x == 7'd594 && y == 7'd375) ||
		(x == 7'd146 && y == 7'd375) || (x == 7'd168 && y == 550) || (x == 452 && y == 7'd272) ||
		(x == 7'd318 && y == 7'd133) || (x == 119 && y == 7'd289) || (x == 204 && y == 7'd361) ||
		(x == 7'd279 && y == 351) || (x == 7'd136 && y == 7'd451) || (x == 7'd362 && y == 7'd531) ||
		(x == 156 && y == 327) || (x == 423 && y == 7'd221) || (x == 279 && y == 7'd108) ||
		(x == 7'd196 && y == 7'd81) || (x == 396 && y == 134) || (x == 7'd632 && y == 7'd391) ||
		(x == 7'd505 && y == 563) || (x == 7'd308 && y == 7'd307) || (x == 7'd402 && y == 7'd505) ||
		(x == 7'd151 && y == 7'd177) || (x == 7'd285 && y == 7'd567) || (x == 7'd100 && y == 634) ||
		(x == 441 && y == 129) || (x == 7'd387 && y == 7'd523) || (x == 7'd271 && y == 7'd216) ||
		(x == 361 && y == 580) || (x == 7'd29 && y == 7'd133) || (x == 7'd503 && y == 7'd619) ||
		(x == 7'd383 && y == 7'd338) || (x == 7'd583 && y == 7'd422) || (x == 157 && y == 159) ||
		(x == 137 && y == 536) || (x == 7'd274 && y == 236) || (x == 269 && y == 7'd116) ||
		(x == 7'd227 && y == 7'd404) || (x == 7'd404 && y == 428) || (x == 7'd222 && y == 625) ||
		(x == 7'd77 && y == 323) || (x == 7'd537 && y == 7'd309) || (x == 7'd410 && y == 7'd48) ||
		(x == 7'd122 && y == 37) || (x == 7'd495 && y == 7) || (x == 7'd71 && y == 7'd130) ||
		(x == 567 && y == 262) || (x == 7'd149 && y == 7'd589) || (x == 7'd634 && y == 7'd141) ||
		(x == 174 && y == 557) || (x == 7'd34 && y == 7'd346) || (x == 7'd630 && y == 7'd345) ||
		(x == 469 && y == 311) || (x == 511 && y == 7'd584) || (x == 351 && y == 7'd264) ||
		(x == 137 && y == 7'd397) || (x == 8 && y == 7'd603) || (x == 7'd449 && y == 7'd227) ||
		(x == 457 && y == 233) || (x == 7'd636 && y == 7'd284) || (x == 222 && y == 7'd14) ||
		(x == 7'd263 && y == 240) || (x == 7'd521 && y == 409) || (x == 7'd545 && y == 7'd628) ||
		(x == 7'd379 && y == 7'd16) || (x == 467 && y == 7'd174) || (x == 7'd540 && y == 7'd354) ||
		(x == 7'd219 && y == 180) || (x == 7'd616 && y == 116) || (x == 7'd18 && y == 3) ||
		(x == 7'd367 && y == 7'd40) || (x == 374 && y == 7'd480) || (x == 509 && y == 204) ||
		(x == 256 && y == 544) || (x == 607 && y == 415) || (x == 7'd241 && y == 7'd216) ||
		(x == 564 && y == 356) || (x == 7'd439 && y == 7'd254) || (x == 7'd87 && y == 7'd122) ||
		(x == 7'd340 && y == 324) || (x == 7'd226 && y == 7'd138) || (x == 7'd343 && y == 7'd105) ||
		(x == 107 && y == 7'd307) || (x == 7'd311 && y == 435) || (x == 532 && y == 7'd600) ||
		(x == 7'd345 && y == 7'd89) || (x == 493 && y == 7'd449) || (x == 519 && y == 491) ||
		(x == 7'd570 && y == 539) || (x == 7'd532 && y == 7'd538) || (x == 7'd375 && y == 86) ||
		(x == 621 && y == 7'd446) || (x == 397 && y == 7'd513) || (x == 7'd366 && y == 456) ||
		(x == 610 && y == 238) || (x == 606 && y == 7'd166) || (x == 289 && y == 422) ||
		(x == 7'd363 && y == 7'd600) || (x == 7'd401 && y == 7'd298) || (x == 7'd167 && y == 7'd397) ||
		(x == 369 && y == 562) || (x == 430 && y == 418) || (x == 7'd343 && y == 7'd371) ||
		(x == 7'd478 && y == 7'd558) || (x == 453 && y == 573) || (x == 141 && y == 329) ||
		(x == 343 && y == 7'd536) || (x == 339 && y == 7'd486) || (x == 7'd523 && y == 7'd467) ||
		(x == 120 && y == 7'd482) || (x == 7'd166 && y == 152) || (x == 466 && y == 499) ||
		(x == 7'd549 && y == 99) || (x == 7'd236 && y == 189) || (x == 7'd522 && y == 7'd62) ||
		(x == 375 && y == 7'd606) || (x == 417 && y == 203) || (x == 34 && y == 7'd339) ||
		(x == 7'd198 && y == 7'd181) || (x == 207 && y == 290) || (x == 608 && y == 7'd600) ||
		(x == 374 && y == 7'd9) || (x == 170 && y == 220) || (x == 160 && y == 598) ||
		(x == 7'd501 && y == 7'd545) || (x == 592 && y == 7'd413) || (x == 7'd22 && y == 437) ||
		(x == 7'd414 && y == 7'd528) || (x == 198 && y == 7'd386) || (x == 466 && y == 7'd266) ||
		(x == 7'd221 && y == 612) || (x == 7'd365 && y == 196) || (x == 626 && y == 317) ||
		(x == 145 && y == 401) || (x == 443 && y == 404) || (x == 587 && y == 190) ||
		(x == 7'd371 && y == 7'd477) || (x == 380 && y == 496) || (x == 166 && y == 192) ||
		(x == 7'd521 && y == 432) || (x == 7'd517 && y == 7'd321) || (x == 609 && y == 608) ||
		(x == 462 && y == 7'd537) || (x == 7'd162 && y == 7'd594) || (x == 7'd118 && y == 335) ||
		(x == 7'd103 && y == 634) || (x == 155 && y == 613) || (x == 440 && y == 621) ||
		(x == 7'd533 && y == 442) || (x == 7'd315 && y == 241) || (x == 7'd286 && y == 556) ||
		(x == 7'd565 && y == 7'd28) || (x == 7'd494 && y == 365) || (x == 515 && y == 7'd530) ||
		(x == 7'd265 && y == 172) || (x == 7'd620 && y == 367) || (x == 339 && y == 7'd600) ||
		(x == 7'd538 && y == 7'd539) || (x == 412 && y == 7'd582) || (x == 528 && y == 7'd319) ||
		(x == 7'd440 && y == 397) || (x == 13 && y == 7'd239) || (x == 302 && y == 214) ||
		(x == 7'd500 && y == 7'd318) || (x == 7'd510 && y == 7'd609) || (x == 7'd564 && y == 416) ||
		(x == 7'd160 && y == 7'd340) || (x == 7'd308 && y == 7'd154) || (x == 7'd551 && y == 7'd145) ||
		(x == 7'd625 && y == 7'd397) || (x == 7'd337 && y == 7'd369) || (x == 7'd0 && y == 332) ||
		(x == 7'd302 && y == 395) || (x == 7'd495 && y == 113) || (x == 331 && y == 478) ||
		(x == 7'd4 && y == 45) || (x == 445 && y == 239) || (x == 7'd448 && y == 46) ||
		(x == 574 && y == 568) || (x == 7'd86 && y == 399) || (x == 7'd249 && y == 7'd137) ||
		(x == 7'd342 && y == 7'd502) || (x == 7'd515 && y == 7'd288) || (x == 7'd188 && y == 7'd449) ||
		(x == 410 && y == 218) || (x == 412 && y == 7'd38) || (x == 7'd338 && y == 7'd191) ||
		(x == 7'd216 && y == 243) || (x == 313 && y == 278) || (x == 185 && y == 219) ||
		(x == 7'd357 && y == 7'd176) || (x == 456 && y == 348) || (x == 313 && y == 7'd392) ||
		(x == 7'd17 && y == 7'd424) || (x == 472 && y == 552) || (x == 606 && y == 317) ||
		(x == 564 && y == 362) || (x == 7'd274 && y == 7'd149) || (x == 322 && y == 229) ||
		(x == 469 && y == 491) || (x == 7'd615 && y == 7'd621) || (x == 333 && y == 358) ||
		(x == 7'd521 && y == 448) || (x == 609 && y == 7'd481) || (x == 7'd577 && y == 7'd230) ||
		(x == 7'd591 && y == 274) || (x == 159 && y == 569) || (x == 7'd80 && y == 296) ||
		(x == 7'd261 && y == 7'd566) || (x == 7'd403 && y == 7'd516) || (x == 7'd379 && y == 7'd334) ||
		(x == 7'd186 && y == 415) || (x == 169 && y == 531) || (x == 7'd354 && y == 545) ||
		(x == 255 && y == 7'd137) || (x == 7'd169 && y == 556) || (x == 7'd122 && y == 160) ||
		(x == 7'd352 && y == 172) || (x == 7'd376 && y == 7'd329) || (x == 7'd65 && y == 7'd248) ||
		(x == 7'd24 && y == 7'd434) || (x == 594 && y == 590) || (x == 7'd556 && y == 145) ||
		(x == 7'd509 && y == 7'd618) || (x == 215 && y == 130) || (x == 530 && y == 577) ||
		(x == 7'd86 && y == 7'd286) || (x == 7'd544 && y == 319) || (x == 7'd600 && y == 499) ||
		(x == 7'd67 && y == 7'd496) || (x == 7'd303 && y == 7'd538) || (x == 486 && y == 250) ||
		(x == 263 && y == 7'd555) || (x == 7'd240 && y == 7'd5) || (x == 547 && y == 7'd64) ||
		(x == 7'd236 && y == 7'd430) || (x == 7'd282 && y == 488) || (x == 555 && y == 585) ||
		(x == 7'd388 && y == 7'd131) || (x == 306 && y == 515) || (x == 452 && y == 7'd170) ||
		(x == 573 && y == 7'd119) || (x == 345 && y == 7'd297) || (x == 7'd543 && y == 7'd449) ||
		(x == 520 && y == 588) || (x == 7'd303 && y == 7) || (x == 7'd388 && y == 308) ||
		(x == 294 && y == 7'd567) || (x == 7'd213 && y == 7'd560) || (x == 510 && y == 7'd239) ||
		(x == 7'd100 && y == 7'd588) || (x == 435 && y == 7'd216) || (x == 559 && y == 7'd144) ||
		(x == 584 && y == 7'd598) || (x == 7'd377 && y == 304) || (x == 7'd317 && y == 7'd505) ||
		(x == 130 && y == 7'd318) || (x == 334 && y == 7'd321) || (x == 421 && y == 289) ||
		(x == 7'd608 && y == 12) || (x == 7'd607 && y == 356) || (x == 7'd214 && y == 534) ||
		(x == 7'd77 && y == 462) || (x == 7'd197 && y == 7'd394) || (x == 458 && y == 7'd399) ||
		(x == 7'd539 && y == 532) || (x == 7'd462 && y == 7'd18) || (x == 7'd562 && y == 317) ||
		(x == 7'd554 && y == 7'd491) || (x == 7'd324 && y == 7'd333) || (x == 7'd532 && y == 7'd195) ||
		(x == 7'd520 && y == 7'd33) || (x == 7'd350 && y == 460) || (x == 7'd511 && y == 532) ||
		(x == 7'd552 && y == 7'd369) || (x == 636 && y == 540) || (x == 358 && y == 7'd219) ||
		(x == 7'd527 && y == 575) || (x == 7'd21 && y == 249) || (x == 138 && y == 7'd227) ||
		(x == 554 && y == 610) || (x == 7'd207 && y == 7'd361) || (x == 267 && y == 326) ||
		(x == 480 && y == 294) || (x == 113 && y == 7'd328) || (x == 7'd466 && y == 193) ||
		(x == 7'd367 && y == 7'd224) || (x == 541 && y == 614) || (x == 7'd402 && y == 7'd152) ||
		(x == 240 && y == 7'd439) || (x == 588 && y == 287) || (x == 360 && y == 7'd319) ||
		(x == 7'd475 && y == 7'd393) || (x == 7'd191 && y == 7'd188) || (x == 242 && y == 149) ||
		(x == 455 && y == 7'd113) || (x == 7'd609 && y == 7'd297) || (x == 233 && y == 7'd430) ||
		(x == 7'd601 && y == 523) || (x == 592 && y == 207) || (x == 7'd188 && y == 7'd134) ||
		(x == 352 && y == 7'd451) || (x == 7'd638 && y == 7'd618) || (x == 276 && y == 535) ||
		(x == 7'd425 && y == 7'd496) || (x == 7'd522 && y == 513) || (x == 7'd454 && y == 7'd165) ||
		(x == 477 && y == 7'd206) || (x == 272 && y == 7'd373) || (x == 156 && y == 7'd126) ||
		(x == 168 && y == 7'd474) || (x == 627 && y == 7'd525) || (x == 7'd365 && y == 227) ||
		(x == 21 && y == 7'd635) || (x == 535 && y == 603) || (x == 7'd326 && y == 7'd73) ||
		(x == 7'd498 && y == 7'd263) || (x == 502 && y == 7'd299) || (x == 7'd615 && y == 569) ||
		(x == 563 && y == 594) || (x == 491 && y == 411) || (x == 403 && y == 7'd225) ||
		(x == 7'd18 && y == 7'd592) || (x == 7'd335 && y == 547) || (x == 223 && y == 133) ||
		(x == 7'd236 && y == 459) || (x == 284 && y == 243) || (x == 7'd351 && y == 7'd337) ||
		(x == 183 && y == 7'd230) || (x == 7'd324 && y == 7'd633) || (x == 356 && y == 639) ||
		(x == 262 && y == 454) || (x == 173 && y == 7'd67) || (x == 124 && y == 7'd274) ||
		(x == 133 && y == 7'd16) || (x == 7'd639 && y == 7'd237) || (x == 192 && y == 181) ||
		(x == 7'd505 && y == 7'd338) || (x == 7'd139 && y == 396) || (x == 7'd539 && y == 7'd389) ||
		(x == 7'd554 && y == 7'd283) || (x == 354 && y == 7'd43) || (x == 7'd141 && y == 7'd472) ||
		(x == 437 && y == 625) || (x == 491 && y == 7'd96) || (x == 7'd588 && y == 170) ||
		(x == 7'd617 && y == 507) || (x == 223 && y == 315) || (x == 264 && y == 382) ||
		(x == 7'd231 && y == 100) || (x == 7'd537 && y == 7'd390) || (x == 7'd223 && y == 7'd295) ||
		(x == 7'd83 && y == 478) || (x == 7'd409 && y == 7'd174) || (x == 572 && y == 7'd636) ||
		(x == 448 && y == 7'd303) || (x == 450 && y == 7'd414) || (x == 7'd233 && y == 7'd301) ||
		(x == 7'd509 && y == 7'd41) || (x == 7'd74 && y == 462) || (x == 156 && y == 302) ||
		(x == 256 && y == 340) || (x == 482 && y == 7'd360) || (x == 637 && y == 7'd194) ||
		(x == 7'd532 && y == 585) || (x == 7'd40 && y == 197) || (x == 7'd144 && y == 7'd321) ||
		(x == 7'd569 && y == 7'd473) || (x == 243 && y == 597) || (x == 7'd63 && y == 7'd521) ||
		(x == 331 && y == 311) || (x == 601 && y == 201) || (x == 228 && y == 570) ||
		(x == 515 && y == 7'd396) || (x == 435 && y == 278) || (x == 7'd472 && y == 7'd243) ||
		(x == 190 && y == 7'd379) || (x == 7'd194 && y == 446) || (x == 367 && y == 330) ||
		(x == 324 && y == 169) || (x == 563 && y == 155) || (x == 7'd614 && y == 7'd286) ||
		(x == 7'd499 && y == 114) || (x == 7'd603 && y == 7'd588) || (x == 394 && y == 7'd379) ||
		(x == 7'd9 && y == 7'd64) || (x == 514 && y == 7'd234) || (x == 556 && y == 7'd183) ||
		(x == 7'd444 && y == 7'd483) || (x == 7'd397 && y == 7'd209) || (x == 126 && y == 7'd360) ||
		(x == 297 && y == 7'd95) || (x == 7'd516 && y == 7'd158) || (x == 408 && y == 402) ||
		(x == 599 && y == 131) || (x == 7'd467 && y == 308) || (x == 7'd288 && y == 502) ||
		(x == 586 && y == 7'd101) || (x == 7'd612 && y == 7'd209) || (x == 616 && y == 7'd197) ||
		(x == 7'd553 && y == 7'd635) || (x == 7'd200 && y == 7'd146) || (x == 403 && y == 239) ||
		(x == 533 && y == 7'd92) || (x == 253 && y == 7'd115) || (x == 7'd592 && y == 7'd112) ||
		(x == 7'd55 && y == 7'd356) || (x == 7'd319 && y == 7'd516) || (x == 7'd246 && y == 7'd585) ||
		(x == 7'd339 && y == 7'd448) || (x == 317 && y == 242) || (x == 7'd624 && y == 7'd191) ||
		(x == 635 && y == 235) || (x == 7'd67 && y == 467) || (x == 7'd375 && y == 553) ||
		(x == 331 && y == 615) || (x == 7'd152 && y == 7'd617) || (x == 7'd27 && y == 400) ||
		(x == 7'd525 && y == 153) || (x == 7'd551 && y == 7'd85) || (x == 609 && y == 7'd565) ||
		(x == 7'd335 && y == 232) || (x == 362 && y == 220) || (x == 7'd189 && y == 7'd602) ||
		(x == 7'd218 && y == 7'd601) || (x == 7'd172 && y == 285) || (x == 323 && y == 7'd286) ||
		(x == 7'd523 && y == 457) || (x == 7'd612 && y == 7'd615) || (x == 595 && y == 7'd360) ||
		(x == 7'd521 && y == 7'd78) || (x == 343 && y == 237) || (x == 171 && y == 344) ||
		(x == 7'd41 && y == 7'd225) || (x == 141 && y == 284) || (x == 453 && y == 339) ||
		(x == 7'd22 && y == 7'd261) || (x == 7'd17 && y == 551) || (x == 7'd429 && y == 210) ||
		(x == 431 && y == 500) || (x == 474 && y == 7'd538) || (x == 292 && y == 132) ||
		(x == 499 && y == 361) || (x == 7'd324 && y == 242) || (x == 7'd320 && y == 7'd305) ||
		(x == 7'd402 && y == 7'd546) || (x == 7'd494 && y == 7'd626) || (x == 525 && y == 7'd550) ||
		(x == 7'd413 && y == 7'd466) || (x == 7'd177 && y == 418) || (x == 536 && y == 187) ||
		(x == 7'd48 && y == 217) || (x == 7'd458 && y == 7'd308) || (x == 374 && y == 7'd400) ||
		(x == 7'd236 && y == 7'd306) || (x == 7'd345 && y == 7) || (x == 7'd267 && y == 7'd245) ||
		(x == 257 && y == 392) || (x == 361 && y == 7'd601) || (x == 271 && y == 7'd0) ||
		(x == 7'd211 && y == 7'd439) || (x == 7'd153 && y == 47) || (x == 7'd15 && y == 117) ||
		(x == 231 && y == 7'd229) || (x == 106 && y == 7'd613) || (x == 638 && y == 7'd424) ||
		(x == 7'd136 && y == 169) || (x == 471 && y == 481) || (x == 204 && y == 203) ||
		(x == 407 && y == 300) || (x == 437 && y == 203) || (x == 7'd563 && y == 431) ||
		(x == 169 && y == 7'd498) || (x == 7'd529 && y == 7'd494) || (x == 7'd306 && y == 310) ||
		(x == 7'd576 && y == 7'd86) || (x == 7'd246 && y == 57) || (x == 7'd241 && y == 7'd575) ||
		(x == 66 && y == 7'd497) || (x == 369 && y == 7'd440) || (x == 294 && y == 444) ||
		(x == 637 && y == 7'd134) || (x == 337 && y == 7'd462) || (x == 7'd230 && y == 7'd309) ||
		(x == 9 && y == 7'd290) || (x == 7'd222 && y == 7'd545) || (x == 7'd332 && y == 7'd348) ||
		(x == 253 && y == 414) || (x == 552 && y == 212) || (x == 7'd378 && y == 579) ||
		(x == 7'd274 && y == 492) || (x == 186 && y == 595) || (x == 400 && y == 569) ||
		(x == 7'd132 && y == 346) || (x == 421 && y == 598) || (x == 159 && y == 462) ||
		(x == 7'd16 && y == 265) || (x == 7'd633 && y == 153) || (x == 636 && y == 451) ||
		(x == 7'd234 && y == 270) || (x == 7'd437 && y == 459) || (x == 7'd618 && y == 275) ||
		(x == 560 && y == 7'd486) || (x == 7'd176 && y == 7'd190) || (x == 7'd496 && y == 200) ||
		(x == 7'd481 && y == 7'd6) || (x == 358 && y == 7'd580) || (x == 7'd53 && y == 469) ||
		(x == 217 && y == 503) || (x == 616 && y == 7'd200) || (x == 573 && y == 577) ||
		(x == 420 && y == 7'd120) || (x == 7'd239 && y == 339) || (x == 7'd496 && y == 7'd284) ||
		(x == 132 && y == 7'd370) || (x == 432 && y == 337) || (x == 7'd297 && y == 390) ||
		(x == 7'd81 && y == 337) || (x == 374 && y == 7'd632) || (x == 434 && y == 536) ||
		(x == 521 && y == 7'd271) || (x == 7'd303 && y == 357) || (x == 7'd544 && y == 425) ||
		(x == 7'd376 && y == 40) || (x == 7'd104 && y == 7'd83) || (x == 7'd81 && y == 384) ||
		(x == 7'd322 && y == 7'd84) || (x == 7'd244 && y == 7'd223) || (x == 102 && y == 7'd262) ||
		(x == 7'd250 && y == 7'd187) || (x == 7'd55 && y == 147) || (x == 568 && y == 322) ||
		(x == 7'd476 && y == 7'd600) || (x == 7'd586 && y == 7'd563) || (x == 7'd62 && y == 7'd225) ||
		(x == 608 && y == 7'd558) || (x == 7'd197 && y == 7'd571) || (x == 7'd423 && y == 629) ||
		(x == 136 && y == 7'd263) || (x == 7'd272 && y == 7'd210) || (x == 7'd141 && y == 559) ||
		(x == 319 && y == 399) || (x == 246 && y == 489) || (x == 7'd16 && y == 360) ||
		(x == 7'd611 && y == 7'd208) || (x == 7'd237 && y == 7'd610) || (x == 7'd503 && y == 293) ||
		(x == 410 && y == 187) || (x == 7'd601 && y == 7'd379) || (x == 7'd371 && y == 7'd624) ||
		(x == 7'd41 && y == 7'd586) || (x == 596 && y == 7'd300) || (x == 602 && y == 182) ||
		(x == 415 && y == 188) || (x == 7'd521 && y == 7'd165) || (x == 7'd303 && y == 7'd8) ||
		(x == 350 && y == 338) || (x == 7'd312 && y == 7'd329) || (x == 7'd367 && y == 7'd567) ||
		(x == 7'd136 && y == 364) || (x == 502 && y == 183) || (x == 151 && y == 483) ||
		(x == 7'd259 && y == 7'd637) || (x == 7'd246 && y == 353) || (x == 552 && y == 351) ||
		(x == 231 && y == 536) || (x == 369 && y == 485) || (x == 7'd168 && y == 187) ||
		(x == 419 && y == 631) || (x == 584 && y == 584) || (x == 7'd225 && y == 580) ||
		(x == 526 && y == 7'd246) || (x == 7'd610 && y == 7'd142) || (x == 7'd256 && y == 344) ||
		(x == 630 && y == 487) || (x == 7'd506 && y == 7'd516) || (x == 172 && y == 392) ||
		(x == 139 && y == 285) || (x == 7'd288 && y == 201) || (x == 7'd497 && y == 532) ||
		(x == 317 && y == 350) || (x == 599 && y == 7'd447) || (x == 7'd576 && y == 7'd141) ||
		(x == 312 && y == 607) || (x == 366 && y == 7'd532) || (x == 7'd283 && y == 483) ||
		(x == 7'd443 && y == 7'd69) || (x == 485 && y == 7'd220) || (x == 7'd490 && y == 566) ||
		(x == 7'd345 && y == 506) || (x == 617 && y == 467) || (x == 450 && y == 190) ||
		(x == 430 && y == 504) || (x == 566 && y == 7'd156) || (x == 7'd608 && y == 7'd550) ||
		(x == 7'd433 && y == 449) || (x == 335 && y == 433) || (x == 434 && y == 298) ||
		(x == 7'd418 && y == 561) || (x == 314 && y == 7'd286) || (x == 7'd227 && y == 7'd437) ||
		(x == 210 && y == 220) || (x == 514 && y == 7'd211) || (x == 7'd155 && y == 231) ||
		(x == 150 && y == 331) || (x == 7'd585 && y == 584) || (x == 7'd548 && y == 408) ||
		(x == 167 && y == 7'd217) || (x == 422 && y == 405) || (x == 340 && y == 363) ||
		(x == 7'd464 && y == 472) || (x == 196 && y == 403) || (x == 7'd562 && y == 565) ||
		(x == 229 && y == 311) || (x == 307 && y == 7'd153) || (x == 7'd580 && y == 7'd546) ||
		(x == 7'd475 && y == 120) || (x == 100 && y == 7'd381) || (x == 7'd581 && y == 446) ||
		(x == 7'd258 && y == 167) || (x == 7'd634 && y == 400) || (x == 292 && y == 354) ||
		(x == 638 && y == 495) || (x == 7'd366 && y == 186) || (x == 28 && y == 7'd129) ||
		(x == 7'd249 && y == 7'd438) || (x == 601 && y == 129) || (x == 168 && y == 488) ||
		(x == 623 && y == 539) || (x == 196 && y == 7'd450) || (x == 7'd488 && y == 7'd209) ||
		(x == 352 && y == 7'd194) || (x == 7'd620 && y == 7'd20) || (x == 7'd492 && y == 7'd633) ||
		(x == 7'd200 && y == 626) || (x == 7'd202 && y == 7'd169) || (x == 7'd449 && y == 410) ||
		(x == 7'd19 && y == 7'd535) || (x == 7'd233 && y == 7'd483) || (x == 7'd163 && y == 7'd471) ||
		(x == 482 && y == 7'd637) || (x == 7'd577 && y == 388) || (x == 7'd603 && y == 7'd272) ||
		(x == 215 && y == 167) || (x == 7'd492 && y == 606) || (x == 7'd85 && y == 168) ||
		(x == 378 && y == 602) || (x == 534 && y == 502) || (x == 7'd440 && y == 570) ||
		(x == 442 && y == 7'd107) || (x == 7'd518 && y == 7'd492) || (x == 575 && y == 7'd214) ||
		(x == 592 && y == 7'd135) || (x == 233 && y == 538) || (x == 7'd198 && y == 7'd508) ||
		(x == 471 && y == 305) || (x == 7'd458 && y == 291) || (x == 7'd556 && y == 7'd200) ||
		(x == 298 && y == 7'd403) || (x == 7'd581 && y == 7'd610) || (x == 448 && y == 480) ||
		(x == 7'd166 && y == 7'd596) || (x == 7'd63 && y == 7'd395) || (x == 7'd45 && y == 241) ||
		(x == 7'd175 && y == 7'd421) || (x == 7'd216 && y == 7'd387) || (x == 71 && y == 7'd263) ||
		(x == 470 && y == 473) || (x == 7'd332 && y == 107) || (x == 7'd455 && y == 7'd495) ||
		(x == 126 && y == 7'd256) || (x == 7'd473 && y == 7'd602) || (x == 284 && y == 583) ||
		(x == 7'd528 && y == 7'd448) || (x == 439 && y == 7'd564) || (x == 219 && y == 7'd453) ||
		(x == 222 && y == 193) || (x == 530 && y == 192) || (x == 7'd629 && y == 13) ||
		(x == 7'd217 && y == 252) || (x == 7'd176 && y == 252) || (x == 7'd556 && y == 7'd583) ||
		(x == 7'd314 && y == 99) || (x == 265 && y == 7'd263) || (x == 7'd340 && y == 7'd563) ||
		(x == 250 && y == 602) || (x == 468 && y == 7'd419) || (x == 7'd238 && y == 454) ||
		(x == 7'd499 && y == 265) || (x == 7'd247 && y == 7'd357) || (x == 226 && y == 7'd383) ||
		(x == 292 && y == 7'd385) || (x == 7'd164 && y == 7'd574) || (x == 7'd576 && y == 7'd448) ||
		(x == 257 && y == 137) || (x == 126 && y == 7'd198) || (x == 7'd291 && y == 7'd404) ||
		(x == 376 && y == 7'd386) || (x == 7'd243 && y == 7'd315) || (x == 169 && y == 380) ||
		(x == 54 && y == 7'd252) || (x == 347 && y == 436) || (x == 7'd538 && y == 636) ||
		(x == 226 && y == 533) || (x == 557 && y == 7'd49) || (x == 227 && y == 7'd441) ||
		(x == 558 && y == 581) || (x == 342 && y == 331) || (x == 7'd550 && y == 7'd158) ||
		(x == 568 && y == 587) || (x == 421 && y == 437) || (x == 519 && y == 7'd185) ||
		(x == 237 && y == 7'd139) || (x == 131 && y == 287) || (x == 593 && y == 7'd595) ||
		(x == 629 && y == 7'd50) || (x == 7'd620 && y == 7'd117) || (x == 172 && y == 592) ||
		(x == 7'd464 && y == 7'd218) || (x == 7'd323 && y == 325) || (x == 7'd93 && y == 195) ||
		(x == 152 && y == 442) || (x == 7'd188 && y == 7'd42) || (x == 7'd536 && y == 498) ||
		(x == 7'd20 && y == 7'd591) || (x == 7'd429 && y == 507) || (x == 7'd427 && y == 7'd84) ||
		(x == 7'd141 && y == 7'd193) || (x == 7'd610 && y == 7'd335) || (x == 122 && y == 39) ||
		(x == 222 && y == 176) || (x == 347 && y == 7'd392) || (x == 7'd460 && y == 7'd556) ||
		(x == 7'd630 && y == 7'd212) || (x == 212 && y == 525) || (x == 7'd41 && y == 268) ||
		(x == 543 && y == 476) || (x == 7'd309 && y == 7'd198) || (x == 7'd504 && y == 7'd96) ||
		(x == 7'd412 && y == 274) || (x == 531 && y == 409) || (x == 7'd61 && y == 418) ||
		(x == 197 && y == 7'd624) || (x == 89 && y == 7'd270) || (x == 235 && y == 531) ||
		(x == 506 && y == 7'd564) || (x == 465 && y == 426) || (x == 233 && y == 322) ||
		(x == 7'd278 && y == 140) || (x == 450 && y == 7'd544) || (x == 7'd156 && y == 7'd271) ||
		(x == 7'd30 && y == 333) || (x == 7'd230 && y == 7'd273) || (x == 7'd442 && y == 7'd253) ||
		(x == 7'd60 && y == 565) || (x == 7'd310 && y == 7'd386) || (x == 157 && y == 401) ||
		(x == 7'd492 && y == 7'd260) || (x == 60 && y == 7'd598) || (x == 7'd474 && y == 7'd143) ||
		(x == 7'd32 && y == 285) || (x == 634 && y == 164) || (x == 7'd40 && y == 240) ||
		(x == 7'd366 && y == 7'd310) || (x == 229 && y == 7'd109) || (x == 516 && y == 7'd166) ||
		(x == 7'd205 && y == 510) || (x == 7'd22 && y == 348) || (x == 7'd178 && y == 7'd258) ||
		(x == 7'd98 && y == 81) || (x == 393 && y == 428) || (x == 7'd193 && y == 7'd475) ||
		(x == 592 && y == 7'd245) || (x == 31 && y == 7'd401) || (x == 447 && y == 163) ||
		(x == 7'd394 && y == 7'd239) || (x == 7'd635 && y == 7'd464) || (x == 562 && y == 626) ||
		(x == 7'd351 && y == 7'd165) || (x == 328 && y == 291) || (x == 7'd359 && y == 7'd426) ||
		(x == 549 && y == 7'd219) || (x == 346 && y == 504) || (x == 467 && y == 7'd454) ||
		(x == 331 && y == 314) || (x == 7'd370 && y == 422) || (x == 300 && y == 485) ||
		(x == 7'd359 && y == 7'd459) || (x == 572 && y == 7'd378) || (x == 110 && y == 7'd374) ||
		(x == 199 && y == 575) || (x == 562 && y == 326) || (x == 7'd184 && y == 522) ||
		(x == 7'd203 && y == 7'd235) || (x == 7'd497 && y == 7'd602) || (x == 7'd571 && y == 180) ||
		(x == 396 && y == 7'd601) || (x == 254 && y == 7'd6) || (x == 7'd31 && y == 7'd580) ||
		(x == 23 && y == 7'd287) || (x == 254 && y == 7'd629) || (x == 577 && y == 7'd599) ||
		(x == 7'd344 && y == 310) || (x == 7'd186 && y == 7'd145) || (x == 7'd101 && y == 216) ||
		(x == 140 && y == 361) || (x == 7'd119 && y == 7'd95) || (x == 238 && y == 7'd87) ||
		(x == 7'd261 && y == 7'd11) || (x == 559 && y == 144) || (x == 7'd209 && y == 7'd224) ||
		(x == 569 && y == 7'd539) || (x == 7'd443 && y == 7'd381) || (x == 7'd299 && y == 7'd376) ||
		(x == 338 && y == 7'd132) || (x == 537 && y == 7'd440) || (x == 43 && y == 7'd286) ||
		(x == 428 && y == 7'd179) || (x == 7'd616 && y == 326) || (x == 7'd579 && y == 7'd633) ||
		(x == 7'd205 && y == 17) || (x == 7'd337 && y == 7'd614) || (x == 595 && y == 7'd66) ||
		(x == 7'd427 && y == 7'd508) || (x == 7'd367 && y == 7'd346) || (x == 455 && y == 7'd16) ||
		(x == 7'd1 && y == 165) || (x == 355 && y == 419) || (x == 7'd405 && y == 7'd307) ||
		(x == 392 && y == 7'd593) || (x == 583 && y == 7'd283) || (x == 362 && y == 292) ||
		(x == 482 && y == 7'd169) || (x == 50 && y == 79) || (x == 7'd619 && y == 502) ||
		(x == 374 && y == 7'd114) || (x == 7'd548 && y == 7'd90) || (x == 428 && y == 339) ||
		(x == 7'd369 && y == 7'd540) || (x == 281 && y == 325) || (x == 7'd151 && y == 7'd160) ||
		(x == 7'd84 && y == 581) || (x == 7'd164 && y == 65) || (x == 7'd211 && y == 7'd513) ||
		(x == 7'd549 && y == 451) || (x == 7'd446 && y == 7'd575) || (x == 7'd185 && y == 416) ||
		(x == 243 && y == 595) || (x == 127 && y == 7'd196) || (x == 165 && y == 176) ||
		(x == 298 && y == 7'd362) || (x == 7'd619 && y == 7'd215) || (x == 7'd626 && y == 7'd445) ||
		(x == 7'd258 && y == 414) || (x == 538 && y == 7'd94) || (x == 155 && y == 7'd50) ||
		(x == 7'd213 && y == 7'd518) || (x == 302 && y == 7'd418) || (x == 7'd580 && y == 581) ||
		(x == 577 && y == 167) || (x == 7'd560 && y == 244) || (x == 7'd594 && y == 7'd555) ||
		(x == 462 && y == 351) || (x == 7'd577 && y == 7'd348) || (x == 381 && y == 413) ||
		(x == 7'd542 && y == 482) || (x == 7'd392 && y == 536) || (x == 7'd375 && y == 574) ||
		(x == 484 && y == 531) || (x == 554 && y == 549) || (x == 591 && y == 410) ||
		(x == 7'd414 && y == 7'd300) || (x == 610 && y == 222) || (x == 7'd497 && y == 11) ||
		(x == 7'd196 && y == 7'd491) || (x == 353 && y == 7'd138) || (x == 7'd533 && y == 464) ||
		(x == 7'd119 && y == 440) || (x == 577 && y == 281) || (x == 7'd457 && y == 7'd614) ||
		(x == 7'd371 && y == 7'd166) || (x == 7'd9 && y == 7'd289) || (x == 110 && y == 7'd281) ||
		(x == 7'd134 && y == 7'd304) || (x == 7'd624 && y == 7'd529) || (x == 299 && y == 211) ||
		(x == 442 && y == 7'd581) || (x == 7'd364 && y == 7'd400) || (x == 7'd370 && y == 7'd442) ||
		(x == 7'd51 && y == 235) || (x == 7'd497 && y == 7'd137) || (x == 409 && y == 7'd32) ||
		(x == 7'd7 && y == 7'd239) || (x == 7'd519 && y == 75) || (x == 302 && y == 308) ||
		(x == 7'd415 && y == 288) || (x == 586 && y == 7'd542) || (x == 265 && y == 7'd152) ||
		(x == 521 && y == 7'd372) || (x == 435 && y == 386) || (x == 403 && y == 602) ||
		(x == 7'd508 && y == 7'd208) || (x == 446 && y == 264) || (x == 229 && y == 7'd333) ||
		(x == 7'd547 && y == 509) || (x == 67 && y == 7'd623) || (x == 7'd532 && y == 7'd524) ||
		(x == 7'd16 && y == 7'd236) || (x == 135 && y == 176) || (x == 7'd115 && y == 7'd509) ||
		(x == 402 && y == 131) || (x == 240 && y == 7'd127) || (x == 7'd307 && y == 7'd363) ||
		(x == 7'd574 && y == 384) || (x == 7'd331 && y == 7'd256) || (x == 7'd212 && y == 151) ||
		(x == 316 && y == 7'd6) || (x == 7'd448 && y == 7'd580) || (x == 7'd520 && y == 393) ||
		(x == 7'd435 && y == 7'd610) || (x == 7'd540 && y == 126) || (x == 230 && y == 7'd280) ||
		(x == 108 && y == 7'd630) || (x == 237 && y == 7'd506) || (x == 7'd373 && y == 7'd320) ||
		(x == 26 && y == 7'd22) || (x == 155 && y == 7'd82) || (x == 627 && y == 193) ||
		(x == 7'd382 && y == 545) || (x == 7'd188 && y == 7'd283) || (x == 629 && y == 7'd300) ||
		(x == 361 && y == 7'd561) || (x == 293 && y == 7'd359) || (x == 7'd90 && y == 7'd560) ||
		(x == 289 && y == 7'd1) || (x == 7'd390 && y == 533) || (x == 197 && y == 142) ||
		(x == 61 && y == 7'd325) || (x == 571 && y == 7'd422) || (x == 7'd565 && y == 7'd329) ||
		(x == 538 && y == 7'd76) || (x == 7'd288 && y == 7'd577) || (x == 249 && y == 238) ||
		(x == 483 && y == 7'd290) || (x == 7'd413 && y == 7'd515) || (x == 595 && y == 443) ||
		(x == 7'd351 && y == 370) || (x == 120 && y == 7'd414) || (x == 242 && y == 7'd34) ||
		(x == 509 && y == 354) || (x == 462 && y == 361) || (x == 233 && y == 281) ||
		(x == 316 && y == 524) || (x == 522 && y == 190) || (x == 634 && y == 171) ||
		(x == 7'd160 && y == 419) || (x == 511 && y == 319) || (x == 7'd161 && y == 7'd460) ||
		(x == 7'd122 && y == 319) || (x == 61 && y == 7'd324) || (x == 7'd406 && y == 7'd633) ||
		(x == 7'd8 && y == 480) || (x == 7'd310 && y == 7'd404) || (x == 7'd521 && y == 7'd243) ||
		(x == 184 && y == 7'd502) || (x == 7'd638 && y == 7'd611) || (x == 7'd486 && y == 124) ||
		(x == 247 && y == 315) || (x == 7'd541 && y == 7'd226) || (x == 613 && y == 453) ||
		(x == 243 && y == 7'd255) || (x == 126 && y == 80) || (x == 591 && y == 281) ||
		(x == 7'd539 && y == 7'd51) || (x == 404 && y == 197) || (x == 7'd382 && y == 7'd460) ||
		(x == 626 && y == 7'd376) || (x == 7'd631 && y == 7'd232) || (x == 610 && y == 258) ||
		(x == 139 && y == 588) || (x == 7'd239 && y == 7'd274) || (x == 7'd41 && y == 7'd270) ||
		(x == 7'd139 && y == 7'd337) || (x == 7'd424 && y == 7'd140) || (x == 7'd570 && y == 7'd450) ||
		(x == 618 && y == 151) || (x == 519 && y == 276) || (x == 605 && y == 7'd117) ||
		(x == 7'd349 && y == 476) || (x == 7'd242 && y == 410) || (x == 7'd570 && y == 366) ||
		(x == 7'd506 && y == 7'd444) || (x == 7'd156 && y == 7'd182) || (x == 7'd177 && y == 565) ||
		(x == 7'd606 && y == 7'd414) || (x == 7'd237 && y == 474) || (x == 7'd549 && y == 7'd630) ||
		(x == 7'd548 && y == 7'd447) || (x == 7'd16 && y == 44) || (x == 249 && y == 633) ||
		(x == 7'd483 && y == 201) || (x == 7'd154 && y == 346) || (x == 7'd12 && y == 7'd245) ||
		(x == 7'd476 && y == 7'd455) || (x == 7'd569 && y == 567) || (x == 152 && y == 7'd133) ||
		(x == 7'd447 && y == 7'd189) || (x == 7'd260 && y == 411) || (x == 514 && y == 7'd37) ||
		(x == 302 && y == 296) || (x == 255 && y == 389) || (x == 618 && y == 7'd32) ||
		(x == 266 && y == 132) || (x == 217 && y == 594) || (x == 7'd616 && y == 405) ||
		(x == 7'd569 && y == 7'd195) || (x == 618 && y == 400) || (x == 617 && y == 7'd506) ||
		(x == 615 && y == 7'd485) || (x == 7'd68 && y == 331) || (x == 7'd46 && y == 38) ||
		(x == 7'd362 && y == 457) || (x == 327 && y == 212) || (x == 7 && y == 7'd527) ||
		(x == 7'd196 && y == 7'd355) || (x == 7'd254 && y == 386) || (x == 616 && y == 7'd557) ||
		(x == 7'd311 && y == 416) || (x == 7'd377 && y == 501) || (x == 504 && y == 7'd101) ||
		(x == 255 && y == 331) || (x == 33 && y == 7'd257) || (x == 566 && y == 7'd333) ||
		(x == 7'd357 && y == 7'd363) || (x == 7'd580 && y == 7'd506) || (x == 110 && y == 7'd343) ||
		(x == 149 && y == 187) || (x == 116 && y == 7'd581) || (x == 7'd614 && y == 100) ||
		(x == 538 && y == 7'd478) || (x == 7'd150 && y == 469) || (x == 532 && y == 7'd378) ||
		(x == 7'd236 && y == 455) || (x == 437 && y == 7'd530) || (x == 535 && y == 7'd516) ||
		(x == 7'd140 && y == 7'd294) || (x == 7'd217 && y == 387) || (x == 7'd22 && y == 7'd285) ||
		(x == 427 && y == 198) || (x == 7'd247 && y == 7'd77) || (x == 7'd237 && y == 556) ||
		(x == 101 && y == 7'd27) || (x == 7'd244 && y == 7'd569) || (x == 7'd143 && y == 570) ||
		(x == 7'd615 && y == 7'd380) || (x == 7'd251 && y == 7'd332) || (x == 161 && y == 345) ||
		(x == 7'd411 && y == 596) || (x == 7'd178 && y == 7'd202) || (x == 499 && y == 7'd116) ||
		(x == 7'd41 && y == 7'd96) || (x == 466 && y == 7'd633) || (x == 7'd383 && y == 71) ||
		(x == 7'd108 && y == 192) || (x == 7'd375 && y == 7'd620) || (x == 7'd415 && y == 7'd464) ||
		(x == 7'd361 && y == 75) || (x == 312 && y == 7'd49) || (x == 596 && y == 7'd271) ||
		(x == 582 && y == 482) || (x == 7'd44 && y == 402) || (x == 302 && y == 387) ||
		(x == 7'd188 && y == 7'd197) || (x == 363 && y == 7'd71) || (x == 7'd274 && y == 1) ||
		(x == 247 && y == 7'd420) || (x == 7'd24 && y == 389) || (x == 7'd498 && y == 7'd164) ||
		(x == 627 && y == 7'd202) || (x == 519 && y == 7'd548) || (x == 7'd240 && y == 7'd542) ||
		(x == 7'd260 && y == 7'd362) || (x == 314 && y == 7'd162) || (x == 267 && y == 7'd415) ||
		(x == 7'd329 && y == 7'd527) || (x == 537 && y == 409) || (x == 151 && y == 311) ||
		(x == 410 && y == 7'd151) || (x == 476 && y == 342) || (x == 386 && y == 7'd339) ||
		(x == 7'd191 && y == 7'd469) || (x == 306 && y == 7'd298) || (x == 7'd398 && y == 7'd552) ||
		(x == 7'd423 && y == 7'd583) || (x == 7'd501 && y == 7'd416) || (x == 7'd542 && y == 7'd449) ||
		(x == 7'd414 && y == 475) || (x == 7'd374 && y == 7'd366) || (x == 7'd577 && y == 7'd373) ||
		(x == 7'd360 && y == 7'd462) || (x == 7'd429 && y == 216) || (x == 148 && y == 7'd363) ||
		(x == 7'd388 && y == 7'd506) || (x == 435 && y == 7'd574) || (x == 82 && y == 7'd430) ||
		(x == 120 && y == 7'd266) || (x == 7'd494 && y == 7'd286) || (x == 7'd507 && y == 7'd447) ||
		(x == 7'd500 && y == 209) || (x == 556 && y == 7'd409) || (x == 7'd388 && y == 7'd565) ||
		(x == 437 && y == 213) || (x == 624 && y == 605) || (x == 371 && y == 7'd610) ||
		(x == 566 && y == 7'd420) || (x == 7'd510 && y == 453) || (x == 487 && y == 7'd550) ||
		(x == 7'd80 && y == 404) || (x == 279 && y == 538) || (x == 7'd137 && y == 7'd602) ||
		(x == 7'd216 && y == 77) || (x == 468 && y == 7'd478) || (x == 476 && y == 7'd581) ||
		(x == 7'd80 && y == 485) || (x == 7'd196 && y == 7'd161) || (x == 7'd322 && y == 47) ||
		(x == 168 && y == 7'd80) || (x == 7'd405 && y == 7'd176) || (x == 7'd393 && y == 370) ||
		(x == 7'd397 && y == 87) || (x == 7'd339 && y == 7'd331) || (x == 203 && y == 7'd388) ||
		(x == 7'd322 && y == 220) || (x == 476 && y == 7'd458) || (x == 353 && y == 216) ||
		(x == 7'd481 && y == 7'd292) || (x == 7'd43 && y == 7'd553) || (x == 165 && y == 7'd181) ||
		(x == 7'd133 && y == 7'd223) || (x == 7'd214 && y == 637) || (x == 7'd573 && y == 7'd528) ||
		(x == 483 && y == 7'd363) || (x == 7'd369 && y == 7'd563) || (x == 557 && y == 7'd147) ||
		(x == 7'd563 && y == 7'd401) || (x == 7'd523 && y == 7'd463) || (x == 7'd299 && y == 12) ||
		(x == 380 && y == 7'd412) || (x == 467 && y == 7'd515) || (x == 534 && y == 520) ||
		(x == 592 && y == 7'd351) || (x == 7'd153 && y == 7'd635) || (x == 417 && y == 7'd541) ||
		(x == 227 && y == 7'd134) || (x == 510 && y == 7'd457) || (x == 7'd113 && y == 7'd252) ||
		(x == 7'd134 && y == 625) || (x == 556 && y == 281) || (x == 7'd72 && y == 263) ||
		(x == 614 && y == 7'd281) || (x == 7'd498 && y == 558) || (x == 7 && y == 7'd366) ||
		(x == 7'd240 && y == 138) || (x == 7'd473 && y == 7'd502) || (x == 7'd439 && y == 312) ||
		(x == 7'd504 && y == 7'd209) || (x == 283 && y == 7'd423) || (x == 7'd345 && y == 208) ||
		(x == 522 && y == 323) || (x == 7'd497 && y == 7'd546) || (x == 7'd250 && y == 606) ||
		(x == 409 && y == 7'd491) || (x == 327 && y == 7'd130) || (x == 459 && y == 7'd618) ||
		(x == 534 && y == 7'd392) || (x == 7'd215 && y == 7'd502) || (x == 254 && y == 141) ||
		(x == 617 && y == 332) || (x == 264 && y == 235) || (x == 226 && y == 7'd272) ||
		(x == 7'd498 && y == 7'd66) || (x == 153 && y == 563) || (x == 7'd623 && y == 7'd599) ||
		(x == 380 && y == 428) || (x == 432 && y == 339) || (x == 558 && y == 320) ||
		(x == 266 && y == 470) || (x == 293 && y == 7'd24) || (x == 7'd488 && y == 605) ||
		(x == 489 && y == 233) || (x == 379 && y == 7'd348) || (x == 153 && y == 7'd329) ||
		(x == 379 && y == 431) || (x == 7'd68 && y == 483) || (x == 7'd372 && y == 533) ||
		(x == 7'd340 && y == 526) || (x == 7'd398 && y == 7'd319) || (x == 7'd364 && y == 97) ||
		(x == 200 && y == 549) || (x == 155 && y == 149) || (x == 7'd471 && y == 7'd505) ||
		(x == 7'd175 && y == 179) || (x == 157 && y == 226) || (x == 7'd281 && y == 419) ||
		(x == 7'd73 && y == 7'd259) || (x == 7'd486 && y == 271) || (x == 7'd354 && y == 599) ||
		(x == 7'd89 && y == 625) || (x == 7'd448 && y == 7'd426) || (x == 635 && y == 374) ||
		(x == 155 && y == 7'd133) || (x == 7'd417 && y == 7'd286) || (x == 7'd194 && y == 7'd458) ||
		(x == 7'd304 && y == 170) || (x == 499 && y == 427) || (x == 7'd55 && y == 194) ||
		(x == 7'd237 && y == 7'd513) || (x == 500 && y == 516) || (x == 7'd588 && y == 7'd351) ||
		(x == 7'd375 && y == 466) || (x == 7'd167 && y == 620) || (x == 7'd637 && y == 528) ||
		(x == 568 && y == 555) || (x == 221 && y == 217) || (x == 453 && y == 7'd385) ||
		(x == 46 && y == 7'd395) || (x == 197 && y == 7'd352) || (x == 479 && y == 7'd1) ||
		(x == 496 && y == 7'd621) || (x == 7'd496 && y == 7'd170) || (x == 331 && y == 326) ||
		(x == 7'd622 && y == 4) || (x == 7'd485 && y == 7'd618) || (x == 7'd636 && y == 7'd593) ||
		(x == 7'd227 && y == 262) || (x == 7'd603 && y == 7'd398) || (x == 171 && y == 302) ||
		(x == 355 && y == 623) || (x == 292 && y == 305) || (x == 7'd360 && y == 7'd432) ||
		(x == 7'd471 && y == 7'd180) || (x == 7'd320 && y == 7'd345) || (x == 7'd59 && y == 562) ||
		(x == 7'd550 && y == 180) || (x == 617 && y == 7'd500) || (x == 7'd406 && y == 7'd125) ||
		(x == 7'd355 && y == 7'd132) || (x == 351 && y == 469) || (x == 448 && y == 526) ||
		(x == 7'd454 && y == 7'd306) || (x == 7'd113 && y == 229) || (x == 6 && y == 7'd195) ||
		(x == 416 && y == 325) || (x == 298 && y == 7'd247) || (x == 7'd193 && y == 7'd115) ||
		(x == 7'd479 && y == 598) || (x == 622 && y == 224) || (x == 7'd239 && y == 7'd322) ||
		(x == 479 && y == 7'd265) || (x == 7'd115 && y == 7'd135) || (x == 608 && y == 7'd566) ||
		(x == 7'd434 && y == 7'd235) || (x == 499 && y == 564) || (x == 7'd296 && y == 7'd14) ||
		(x == 7'd422 && y == 184) || (x == 554 && y == 7'd395) || (x == 113 && y == 7'd509) ||
		(x == 7'd435 && y == 593) || (x == 230 && y == 386) || (x == 7'd377 && y == 7'd208) ||
		(x == 504 && y == 431) || (x == 319 && y == 288) || (x == 7'd6 && y == 7'd428) ||
		(x == 75 && y == 17) || (x == 280 && y == 7'd440) || (x == 7'd406 && y == 249) ||
		(x == 7'd173 && y == 423) || (x == 414 && y == 7'd392) || (x == 235 && y == 7'd529) ||
		(x == 318 && y == 454) || (x == 7'd344 && y == 7'd247) || (x == 7'd88 && y == 30) ||
		(x == 7'd74 && y == 364) || (x == 7'd608 && y == 7'd583) || (x == 7'd395 && y == 7'd405) ||
		(x == 7'd359 && y == 7'd507) || (x == 7'd603 && y == 7'd419) || (x == 7'd288 && y == 7'd209) ||
		(x == 7'd41 && y == 7'd634) || (x == 7'd509 && y == 592) || (x == 7'd377 && y == 7'd60) ||
		(x == 291 && y == 7'd570) || (x == 473 && y == 403) || (x == 89 && y == 7'd245) ||
		(x == 7'd108 && y == 7'd227) || (x == 7'd191 && y == 7'd263) || (x == 7'd402 && y == 7'd548) ||
		(x == 527 && y == 354) || (x == 7'd176 && y == 7'd508) || (x == 255 && y == 7'd595) ||
		(x == 7'd413 && y == 7'd196) || (x == 7'd574 && y == 114) || (x == 352 && y == 7'd169) ||
		(x == 557 && y == 295) || (x == 7'd637 && y == 7'd589) || (x == 7'd167 && y == 7'd1) ||
		(x == 7'd143 && y == 492) || (x == 537 && y == 481) || (x == 7'd461 && y == 489) ||
		(x == 227 && y == 7'd17) || (x == 7'd62 && y == 460) || (x == 339 && y == 352) ||
		(x == 7'd539 && y == 7'd491) || (x == 7'd10 && y == 7'd417) || (x == 421 && y == 615) ||
		(x == 438 && y == 231) || (x == 7'd33 && y == 180) || (x == 87 && y == 7'd372) ||
		(x == 7'd635 && y == 7'd269) || (x == 7'd363 && y == 251) || (x == 30 && y == 7'd223) ||
		(x == 7'd324 && y == 7'd164) || (x == 256 && y == 324) || (x == 7'd451 && y == 7'd419) ||
		(x == 7'd9 && y == 7'd291) || (x == 7'd606 && y == 514) || (x == 7'd579 && y == 465) ||
		(x == 7'd120 && y == 7'd506) || (x == 540 && y == 7'd140) || (x == 7'd321 && y == 313) ||
		(x == 7'd407 && y == 7'd174) || (x == 7'd354 && y == 7'd622) || (x == 7'd518 && y == 307) ||
		(x == 242 && y == 267) || (x == 167 && y == 372) || (x == 7'd273 && y == 7'd164) ||
		(x == 7'd9 && y == 7'd314) || (x == 7'd506 && y == 251) || (x == 7'd530 && y == 7'd85) ||
		(x == 390 && y == 137) || (x == 7'd241 && y == 7'd413) || (x == 7'd613 && y == 603) ||
		(x == 7'd278 && y == 438) || (x == 7'd624 && y == 7'd636) || (x == 7'd392 && y == 7'd554) ||
		(x == 268 && y == 272) || (x == 7'd453 && y == 7'd262) || (x == 430 && y == 7'd458) ||
		(x == 7'd59 && y == 368) || (x == 258 && y == 594) || (x == 7'd412 && y == 7'd633) ||
		(x == 137 && y == 604) || (x == 7'd469 && y == 7'd261) || (x == 7'd624 && y == 414) ||
		(x == 378 && y == 630) || (x == 10 && y == 7'd346) || (x == 7'd290 && y == 7'd384) ||
		(x == 444 && y == 7'd295) || (x == 231 && y == 7'd448) || (x == 7'd507 && y == 7'd361) ||
		(x == 71 && y == 7'd17) || (x == 552 && y == 7'd25) || (x == 7'd5 && y == 7'd235) ||
		(x == 530 && y == 354) || (x == 284 && y == 336) || (x == 7'd546 && y == 577) ||
		(x == 26 && y == 13) || (x == 500 && y == 7'd532) || (x == 7'd162 && y == 409) ||
		(x == 7'd230 && y == 7'd121) || (x == 390 && y == 7'd24) || (x == 7'd525 && y == 7'd113) ||
		(x == 631 && y == 338) || (x == 7'd87 && y == 142) || (x == 271 && y == 7'd183) ||
		(x == 475 && y == 7'd209) || (x == 376 && y == 552) || (x == 7'd447 && y == 638) ||
		(x == 7'd370 && y == 68) || (x == 474 && y == 620) || (x == 7'd266 && y == 7'd66) ||
		(x == 522 && y == 7'd623) || (x == 186 && y == 635) || (x == 7'd474 && y == 95) ||
		(x == 7'd480 && y == 7'd264) || (x == 191 && y == 7'd161) || (x == 7'd39 && y == 7'd144) ||
		(x == 7'd4 && y == 7'd360) || (x == 404 && y == 7'd161) || (x == 7'd618 && y == 7'd560) ||
		(x == 7'd616 && y == 7'd170) || (x == 593 && y == 7'd488) || (x == 7'd175 && y == 7'd591) ||
		(x == 7'd265 && y == 7'd299) || (x == 188 && y == 7'd556) || (x == 449 && y == 7'd526) ||
		(x == 7'd105 && y == 7'd338) || (x == 7'd457 && y == 466) || (x == 212 && y == 7'd53) ||
		(x == 7'd572 && y == 7'd112) || (x == 344 && y == 524) || (x == 7'd314 && y == 347) ||
		(x == 7'd592 && y == 415) || (x == 7'd361 && y == 7'd129) || (x == 266 && y == 7'd382) ||
		(x == 7'd576 && y == 229) || (x == 625 && y == 7'd444) || (x == 7'd270 && y == 7'd512) ||
		(x == 7'd553 && y == 230) || (x == 512 && y == 7'd327) || (x == 7'd179 && y == 375) ||
		(x == 7'd631 && y == 7'd204) || (x == 7'd417 && y == 361) || (x == 7'd74 && y == 210) ||
		(x == 610 && y == 7'd404) || (x == 69 && y == 7'd177) || (x == 153 && y == 7'd382) ||
		(x == 556 && y == 374) || (x == 507 && y == 474) || (x == 7'd306 && y == 335) ||
		(x == 7'd253 && y == 7'd128) || (x == 7'd616 && y == 7'd357) || (x == 548 && y == 313) ||
		(x == 7'd628 && y == 7'd7) || (x == 187 && y == 357) || (x == 637 && y == 7'd113) ||
		(x == 7'd211 && y == 267) || (x == 7'd223 && y == 446) || (x == 552 && y == 7'd253) ||
		(x == 7'd497 && y == 62) || (x == 7'd276 && y == 7'd525) || (x == 7'd431 && y == 7'd140) ||
		(x == 7'd433 && y == 588) || (x == 7'd116 && y == 268) || (x == 7'd261 && y == 7'd7) ||
		(x == 7'd360 && y == 7'd583) || (x == 7'd583 && y == 578) || (x == 439 && y == 7'd361) ||
		(x == 7'd387 && y == 7'd159) || (x == 7'd204 && y == 7'd225) || (x == 7'd57 && y == 537) ||
		(x == 7'd388 && y == 581) || (x == 7'd230 && y == 637) || (x == 7'd266 && y == 7'd404) ||
		(x == 345 && y == 7'd327) || (x == 7'd574 && y == 375) || (x == 235 && y == 292) ||
		(x == 7'd57 && y == 185) || (x == 327 && y == 154) || (x == 530 && y == 340) ||
		(x == 225 && y == 7'd37) || (x == 7'd614 && y == 165) || (x == 194 && y == 7'd483) ||
		(x == 7'd413 && y == 7'd325) || (x == 7'd19 && y == 240) || (x == 7'd466 && y == 7'd628) ||
		(x == 381 && y == 7'd425) || (x == 7'd473 && y == 7'd37) || (x == 7'd530 && y == 7'd161) ||
		(x == 7'd270 && y == 7'd468) || (x == 354 && y == 287) || (x == 626 && y == 545) ||
		(x == 7'd64 && y == 161) || (x == 7'd399 && y == 614) || (x == 7'd581 && y == 7'd204) ||
		(x == 7'd59 && y == 7'd506) || (x == 7'd516 && y == 7'd233) || (x == 7'd69 && y == 554) ||
		(x == 404 && y == 401) || (x == 7'd270 && y == 7'd528) || (x == 575 && y == 7'd512) ||
		(x == 553 && y == 7'd229) || (x == 7'd103 && y == 7'd588) || (x == 7'd613 && y == 7'd275) ||
		(x == 409 && y == 519) || (x == 301 && y == 511) || (x == 7'd76 && y == 7'd83) ||
		(x == 7'd475 && y == 7'd455) || (x == 7'd66 && y == 7'd186) || (x == 147 && y == 270) ||
		(x == 7'd260 && y == 411) || (x == 45 && y == 7'd134) || (x == 7'd433 && y == 571) ||
		(x == 572 && y == 7'd595) || (x == 7'd328 && y == 7'd294) || (x == 7'd277 && y == 7'd263) ||
		(x == 7'd293 && y == 584) || (x == 7'd226 && y == 6) || (x == 273 && y == 205) ||
		(x == 7'd494 && y == 7'd560) || (x == 7'd557 && y == 7'd251) || (x == 7'd126 && y == 315) ||
		(x == 144 && y == 632) || (x == 7'd485 && y == 7'd295) || (x == 153 && y == 7'd41) ||
		(x == 415 && y == 7'd225) || (x == 313 && y == 193) || (x == 436 && y == 154) ||
		(x == 415 && y == 482) || (x == 587 && y == 542) || (x == 7'd318 && y == 7'd139) ||
		(x == 222 && y == 239) || (x == 7'd405 && y == 7'd247) || (x == 7'd469 && y == 402) ||
		(x == 7'd510 && y == 7'd371) || (x == 7'd274 && y == 7'd58) || (x == 7'd88 && y == 530) ||
		(x == 7'd83 && y == 7'd66) || (x == 7'd253 && y == 56) || (x == 7'd29 && y == 372) ||
		(x == 164 && y == 7'd602) || (x == 552 && y == 161) || (x == 7'd335 && y == 330) ||
		(x == 391 && y == 7'd418) || (x == 7'd37 && y == 7'd375) || (x == 7'd628 && y == 7'd65) ||
		(x == 277 && y == 451) || (x == 7'd118 && y == 328) || (x == 7'd335 && y == 7'd624) ||
		(x == 428 && y == 289) || (x == 640 && y == 433) || (x == 7'd243 && y == 435) ||
		(x == 284 && y == 411) || (x == 7'd380 && y == 7'd427) || (x == 7'd216 && y == 7'd473) ||
		(x == 570 && y == 7'd428) || (x == 7'd476 && y == 553) || (x == 297 && y == 271) ||
		(x == 443 && y == 7'd562) || (x == 552 && y == 354) || (x == 7'd509 && y == 7'd411) ||
		(x == 7'd239 && y == 7'd288) || (x == 479 && y == 7'd310) || (x == 7'd261 && y == 7'd455) ||
		(x == 181 && y == 7'd140) || (x == 90 && y == 7'd542) || (x == 351 && y == 215) ||
		(x == 7'd460 && y == 7'd0) || (x == 7'd567 && y == 7'd257) || (x == 7'd216 && y == 50) ||
		(x == 7'd233 && y == 7'd377) || (x == 7'd382 && y == 7'd356) || (x == 7'd306 && y == 218) ||
		(x == 7'd491 && y == 7'd1) || (x == 7'd198 && y == 7'd183) || (x == 453 && y == 7'd451) ||
		(x == 7'd364 && y == 7'd605) || (x == 7'd330 && y == 371) || (x == 7'd629 && y == 147) ||
		(x == 7'd507 && y == 14) || (x == 638 && y == 157) || (x == 65 && y == 119) ||
		(x == 7'd26 && y == 372) || (x == 568 && y == 234) || (x == 7'd593 && y == 7'd607) ||
		(x == 7'd397 && y == 37) || (x == 7'd5 && y == 7'd286) || (x == 135 && y == 588) ||
		(x == 457 && y == 7'd329) || (x == 7'd541 && y == 7'd171) || (x == 632 && y == 7'd305) ||
		(x == 7'd449 && y == 392) || (x == 7'd90 && y == 7'd583) || (x == 487 && y == 157) ||
		(x == 456 && y == 7'd308) || (x == 7'd416 && y == 219) || (x == 7'd148 && y == 7'd280) ||
		(x == 7'd236 && y == 7'd370) || (x == 446 && y == 613) || (x == 524 && y == 7'd372) ||
		(x == 7'd507 && y == 7'd438) || (x == 279 && y == 7'd525) || (x == 599 && y == 7'd441) ||
		(x == 7'd571 && y == 634) || (x == 7'd541 && y == 7'd322) || (x == 7'd395 && y == 7'd19) ||
		(x == 7'd302 && y == 7'd394) || (x == 7'd499 && y == 7'd54) || (x == 7'd273 && y == 7'd549) ||
		(x == 7'd451 && y == 7'd353) || (x == 7'd179 && y == 7'd389) || (x == 7'd549 && y == 7'd217) ||
		(x == 280 && y == 315) || (x == 7'd45 && y == 7'd141) || (x == 7'd305 && y == 403) ||
		(x == 157 && y == 187) || (x == 414 && y == 7'd444) || (x == 531 && y == 7'd51) ||
		(x == 7'd163 && y == 7'd66) || (x == 7'd504 && y == 7'd380) || (x == 7'd117 && y == 563) ||
		(x == 529 && y == 238) || (x == 7'd50 && y == 7'd204) || (x == 7'd321 && y == 7'd45) ||
		(x == 271 && y == 617) || (x == 7'd339 && y == 7'd572) || (x == 321 && y == 7'd441) ||
		(x == 269 && y == 413) || (x == 159 && y == 262) || (x == 7'd516 && y == 7'd327) ||
		(x == 497 && y == 615) || (x == 7'd520 && y == 409) || (x == 355 && y == 435) ||
		(x == 393 && y == 303) || (x == 302 && y == 499) || (x == 396 && y == 7'd498) ||
		(x == 7'd106 && y == 7'd595) || (x == 7'd267 && y == 7'd444) || (x == 550 && y == 7'd71) ||
		(x == 7'd5 && y == 7'd92) || (x == 7'd8 && y == 533) || (x == 445 && y == 249) ||
		(x == 155 && y == 7'd77) || (x == 7'd377 && y == 7'd186) || (x == 7'd3 && y == 554) ||
		(x == 7'd455 && y == 271) || (x == 280 && y == 592) || (x == 7'd467 && y == 7'd69) ||
		(x == 7'd407 && y == 389) || (x == 7'd570 && y == 7'd341) || (x == 7'd200 && y == 346) ||
		(x == 7'd578 && y == 92) || (x == 7'd135 && y == 7'd56) || (x == 7'd309 && y == 7'd275) ||
		(x == 133 && y == 341) || (x == 7'd198 && y == 56) || (x == 7'd478 && y == 8) ||
		(x == 632 && y == 7'd368) || (x == 7'd267 && y == 7'd144) || (x == 239 && y == 7'd94) ||
		(x == 623 && y == 7'd406) || (x == 7'd231 && y == 7'd171) || (x == 506 && y == 371) ||
		(x == 7'd584 && y == 7'd460) || (x == 7'd351 && y == 7'd164) || (x == 7'd13 && y == 203) ||
		(x == 298 && y == 7'd513) || (x == 559 && y == 7'd429) || (x == 7'd147 && y == 429) ||
		(x == 7'd490 && y == 152) || (x == 7'd29 && y == 7'd269) || (x == 129 && y == 7'd588) ||
		(x == 162 && y == 7'd192) || (x == 7'd598 && y == 7'd536) || (x == 7'd314 && y == 420) ||
		(x == 569 && y == 7'd374) || (x == 186 && y == 7'd231) || (x == 7'd555 && y == 7'd238) ||
		(x == 378 && y == 7'd146) || (x == 282 && y == 7'd200) || (x == 558 && y == 7'd331) ||
		(x == 615 && y == 7'd443) || (x == 175 && y == 480) || (x == 7'd326 && y == 14) ||
		(x == 451 && y == 602) || (x == 7'd376 && y == 7'd355) || (x == 469 && y == 169) ||
		(x == 238 && y == 573) || (x == 637 && y == 7'd505) || (x == 134 && y == 7'd404) ||
		(x == 7'd546 && y == 465) || (x == 467 && y == 7'd316) || (x == 537 && y == 596) ||
		(x == 7'd581 && y == 7'd165) || (x == 154 && y == 489) || (x == 501 && y == 7'd444) ||
		(x == 7'd5 && y == 7'd578) || (x == 7'd134 && y == 7'd543) || (x == 7'd147 && y == 7'd506) ||
		(x == 544 && y == 576) || (x == 361 && y == 7'd138) || (x == 196 && y == 129) ||
		(x == 297 && y == 338) || (x == 327 && y == 518) || (x == 7'd93 && y == 130) ||
		(x == 256 && y == 436) || (x == 563 && y == 7'd492) || (x == 7'd631 && y == 7'd469) ||
		(x == 565 && y == 165) || (x == 7'd100 && y == 7'd507) || (x == 7'd284 && y == 461) ||
		(x == 350 && y == 7'd47) || (x == 43 && y == 7'd230) || (x == 163 && y == 290) ||
		(x == 166 && y == 216) || (x == 7'd180 && y == 7'd16) || (x == 572 && y == 7'd303) ||
		(x == 448 && y == 7'd355) || (x == 7'd11 && y == 7'd446) || (x == 7'd373 && y == 7'd183) ||
		(x == 525 && y == 544) || (x == 7'd615 && y == 7'd505) || (x == 510 && y == 7'd305) ||
		(x == 223 && y == 637) || (x == 7'd248 && y == 7'd249) || (x == 7'd259 && y == 571) ||
		(x == 129 && y == 7'd636) || (x == 608 && y == 168) || (x == 339 && y == 487) ||
		(x == 342 && y == 368) || (x == 7'd157 && y == 7'd456) || (x == 7'd243 && y == 192) ||
		(x == 237 && y == 247) || (x == 7'd55 && y == 7'd623) || (x == 7'd634 && y == 7'd544) ||
		(x == 506 && y == 7'd468) || (x == 124 && y == 7'd55) || (x == 7'd577 && y == 7'd113) ||
		(x == 311 && y == 418) || (x == 213 && y == 7'd63) || (x == 139 && y == 7'd588) ||
		(x == 421 && y == 7'd116) || (x == 7'd386 && y == 144) || (x == 161 && y == 7'd34) ||
		(x == 7'd498 && y == 214) || (x == 7'd627 && y == 7'd239) || (x == 418 && y == 221) ||
		(x == 6 && y == 7'd183) || (x == 7'd474 && y == 7'd627) || (x == 614 && y == 7'd10) ||
		(x == 7'd56 && y == 225) || (x == 7'd548 && y == 274) || (x == 7'd540 && y == 319) ||
		(x == 461 && y == 7'd68) || (x == 260 && y == 7'd325) || (x == 7'd195 && y == 7'd265) ||
		(x == 7'd267 && y == 434) || (x == 432 && y == 7'd64) || (x == 7'd584 && y == 7'd400) ||
		(x == 423 && y == 7'd416) || (x == 574 && y == 7'd475) || (x == 7'd241 && y == 30) ||
		(x == 7'd121 && y == 7'd635) || (x == 182 && y == 7'd493) || (x == 452 && y == 7'd388) ||
		(x == 305 && y == 181) || (x == 7'd551 && y == 624) || (x == 7'd248 && y == 7'd381) ||
		(x == 7'd635 && y == 7'd340) || (x == 499 && y == 239) || (x == 485 && y == 591) ||
		(x == 402 && y == 257) || (x == 7'd34 && y == 570) || (x == 7'd30 && y == 7'd197) ||
		(x == 7'd217 && y == 623) || (x == 490 && y == 7'd446) || (x == 7'd443 && y == 7'd218) ||
		(x == 7'd598 && y == 1) || (x == 7'd134 && y == 7'd91) || (x == 206 && y == 160) ||
		(x == 20 && y == 7'd182) || (x == 296 && y == 7'd476) || (x == 7'd208 && y == 7'd126) ||
		(x == 7'd132 && y == 24) || (x == 7'd396 && y == 7'd463) || (x == 7'd431 && y == 7'd283) ||
		(x == 7'd143 && y == 7'd535) || (x == 172 && y == 533) || (x == 7'd112 && y == 7'd274) ||
		(x == 606 && y == 7'd206) || (x == 207 && y == 283) || (x == 7'd541 && y == 288) ||
		(x == 7'd252 && y == 7'd309) || (x == 7'd129 && y == 615) || (x == 7'd518 && y == 7'd332) ||
		(x == 7'd522 && y == 7'd466) || (x == 585 && y == 7'd535) || (x == 269 && y == 482) ||
		(x == 7'd136 && y == 7'd108) || (x == 252 && y == 7'd398) || (x == 7'd163 && y == 7'd348) ||
		(x == 630 && y == 7'd277) || (x == 299 && y == 7'd280) || (x == 593 && y == 7'd449) ||
		(x == 7'd238 && y == 7'd342) || (x == 187 && y == 7'd522) || (x == 7'd524 && y == 7'd208) ||
		(x == 530 && y == 338) || (x == 7'd418 && y == 375) || (x == 310 && y == 7'd19) ||
		(x == 7'd521 && y == 7'd129) || (x == 179 && y == 7'd428) || (x == 458 && y == 381) ||
		(x == 317 && y == 7'd299) || (x == 406 && y == 409) || (x == 240 && y == 311) ||
		(x == 7'd205 && y == 7'd601) || (x == 7'd399 && y == 467) || (x == 7'd636 && y == 7'd632) ||
		(x == 7'd296 && y == 618) || (x == 418 && y == 274) || (x == 597 && y == 139) ||
		(x == 7'd271 && y == 7'd256) || (x == 174 && y == 7'd324) || (x == 7'd583 && y == 130) ||
		(x == 344 && y == 547) || (x == 7'd457 && y == 7'd254) || (x == 510 && y == 7'd76) ||
		(x == 7'd98 && y == 7'd552) || (x == 166 && y == 322) || (x == 7'd460 && y == 7'd130) ||
		(x == 386 && y == 612) || (x == 7'd186 && y == 576) || (x == 33 && y == 7'd211) ||
		(x == 386 && y == 7'd451) || (x == 7'd15 && y == 421) || (x == 477 && y == 7'd500) ||
		(x == 7'd510 && y == 7'd433) || (x == 354 && y == 7'd224) || (x == 7'd510 && y == 7'd435) ||
		(x == 7'd272 && y == 141) || (x == 297 && y == 7'd627) || (x == 587 && y == 7'd546) ||
		(x == 178 && y == 199) || (x == 563 && y == 7'd444) || (x == 7'd392 && y == 7'd491) ||
		(x == 7'd189 && y == 7'd46) || (x == 406 && y == 335) || (x == 473 && y == 330) ||
		(x == 7'd505 && y == 455) || (x == 640 && y == 188) || (x == 7'd114 && y == 607) ||
		(x == 7'd608 && y == 7'd431) || (x == 7'd363 && y == 7'd515) || (x == 7'd532 && y == 7'd521) ||
		(x == 7'd550 && y == 7'd587) || (x == 7'd571 && y == 7'd259) || (x == 460 && y == 7'd35) ||
		(x == 7'd551 && y == 7'd248) || (x == 7'd191 && y == 349) || (x == 7'd480 && y == 7'd382) ||
		(x == 355 && y == 584) || (x == 26 && y == 7'd407) || (x == 7'd15 && y == 7'd423) ||
		(x == 359 && y == 7'd127) || (x == 7'd452 && y == 436) || (x == 7'd594 && y == 7'd582) ||
		(x == 424 && y == 243) || (x == 7'd412 && y == 7'd82) || (x == 7'd578 && y == 7'd503) ||
		(x == 7'd231 && y == 99) || (x == 7'd235 && y == 7'd115) || (x == 259 && y == 7'd147) ||
		(x == 439 && y == 7'd32) || (x == 7'd281 && y == 7'd305) || (x == 63 && y == 7'd505) ||
		(x == 7'd275 && y == 1) || (x == 532 && y == 221) || (x == 7'd205 && y == 413) ||
		(x == 239 && y == 7'd263) || (x == 7'd552 && y == 7'd216) || (x == 7'd297 && y == 428) ||
		(x == 7'd399 && y == 433) || (x == 129 && y == 7'd531) || (x == 7'd526 && y == 7'd630) ||
		(x == 565 && y == 7'd175) || (x == 7'd469 && y == 353) || (x == 543 && y == 474) ||
		(x == 612 && y == 511) || (x == 40 && y == 7'd445) || (x == 7'd380 && y == 273) ||
		(x == 7'd65 && y == 7'd473) || (x == 7'd105 && y == 7'd354) || (x == 7'd228 && y == 7'd594) ||
		(x == 7'd161 && y == 7'd549) || (x == 141 && y == 520) || (x == 7'd521 && y == 7'd400) ||
		(x == 557 && y == 502) || (x == 146 && y == 380) || (x == 7'd354 && y == 7'd164) ||
		(x == 381 && y == 7'd311) || (x == 7'd444 && y == 7'd370) || (x == 7'd521 && y == 63) ||
		(x == 201 && y == 625) || (x == 7'd417 && y == 7'd604) || (x == 584 && y == 166) ||
		(x == 7'd253 && y == 7'd208) || (x == 7'd286 && y == 125) || (x == 7'd365 && y == 0) ||
		(x == 7'd453 && y == 393) || (x == 7'd88 && y == 467) || (x == 491 && y == 7'd588) ||
		(x == 7'd254 && y == 7'd559) || (x == 7'd17 && y == 633) || (x == 7'd12 && y == 520) ||
		(x == 28 && y == 7'd565) || (x == 7'd404 && y == 7'd380) || (x == 7'd203 && y == 478) ||
		(x == 7'd443 && y == 7'd472) || (x == 7'd435 && y == 7'd223) || (x == 275 && y == 7'd312) ||
		(x == 7'd297 && y == 7'd516) || (x == 525 && y == 433) || (x == 335 && y == 7'd284) ||
		(x == 7'd610 && y == 7'd231) || (x == 7'd590 && y == 7'd111) || (x == 7'd590 && y == 7'd327) ||
		(x == 7'd332 && y == 7'd90) || (x == 473 && y == 235) || (x == 320 && y == 508) ||
		(x == 511 && y == 7'd422) || (x == 7'd537 && y == 182) || (x == 316 && y == 151) ||
		(x == 545 && y == 7'd378) || (x == 153 && y == 7'd503) || (x == 7'd111 && y == 7'd437) ||
		(x == 321 && y == 333) || (x == 7'd32 && y == 337) || (x == 7'd373 && y == 7'd440) ||
		(x == 7'd350 && y == 7'd53) || (x == 7'd222 && y == 7'd160) || (x == 7'd327 && y == 7'd396) ||
		(x == 7'd519 && y == 7'd619) || (x == 560 && y == 7'd283) || (x == 7'd151 && y == 28) ||
		(x == 622 && y == 411) || (x == 7'd458 && y == 182) || (x == 7'd355 && y == 7'd549) ||
		(x == 7'd148 && y == 7'd290) || (x == 7'd448 && y == 7'd506) || (x == 7'd558 && y == 7'd233) ||
		(x == 454 && y == 360) || (x == 52 && y == 7'd361) || (x == 7'd275 && y == 7'd237) ||
		(x == 636 && y == 7'd420) || (x == 412 && y == 627) || (x == 155 && y == 7'd550) ||
		(x == 324 && y == 7'd352) || (x == 479 && y == 7'd244) || (x == 7'd196 && y == 7'd498) ||
		(x == 7'd171 && y == 7'd583) || (x == 7'd331 && y == 424) || (x == 625 && y == 318) ||
		(x == 7'd391 && y == 34) || (x == 7'd37 && y == 7'd163) || (x == 7'd431 && y == 373) ||
		(x == 274 && y == 266) || (x == 7'd518 && y == 7'd24) || (x == 7'd594 && y == 7'd187) ||
		(x == 526 && y == 321) || (x == 456 && y == 7'd25) || (x == 7'd86 && y == 323) ||
		(x == 7'd423 && y == 533) || (x == 7'd75 && y == 425) || (x == 7'd438 && y == 225) ||
		(x == 7'd575 && y == 7'd301) || (x == 7'd118 && y == 221) || (x == 7'd316 && y == 7'd599) ||
		(x == 186 && y == 7'd277) || (x == 7'd225 && y == 7'd361) || (x == 7'd584 && y == 630) ||
		(x == 548 && y == 340) || (x == 625 && y == 343) || (x == 218 && y == 7'd235) ||
		(x == 451 && y == 580) || (x == 7'd624 && y == 230) || (x == 7'd338 && y == 7'd563) ||
		(x == 7'd337 && y == 7'd128) || (x == 511 && y == 7'd214) || (x == 7'd398 && y == 358) ||
		(x == 459 && y == 307) || (x == 7'd387 && y == 7'd133) || (x == 197 && y == 485) ||
		(x == 162 && y == 155) || (x == 293 && y == 407) || (x == 7'd348 && y == 359) ||
		(x == 4 && y == 10) || (x == 7'd319 && y == 156) || (x == 7'd515 && y == 7'd325) ||
		(x == 7'd214 && y == 7'd608) || (x == 346 && y == 241) || (x == 8 && y == 7'd152) ||
		(x == 7'd160 && y == 465) || (x == 21 && y == 7'd302) || (x == 98 && y == 17) ||
		(x == 572 && y == 369) || (x == 410 && y == 503) || (x == 7'd441 && y == 435) ||
		(x == 276 && y == 7'd584) || (x == 7'd575 && y == 386) || (x == 7'd8 && y == 34) ||
		(x == 7'd42 && y == 7'd118) || (x == 7'd600 && y == 224) || (x == 7'd229 && y == 123) ||
		(x == 7'd378 && y == 7'd387) || (x == 7'd80 && y == 7'd215) || (x == 7'd75 && y == 620) ||
		(x == 7'd93 && y == 301) || (x == 161 && y == 399) || (x == 131 && y == 7'd445) ||
		(x == 7'd242 && y == 7'd447) || (x == 268 && y == 553) || (x == 370 && y == 610) ||
		(x == 83 && y == 7'd174) || (x == 7'd350 && y == 108) || (x == 7'd482 && y == 7'd393) ||
		(x == 58 && y == 7'd16) || (x == 7'd625 && y == 254) || (x == 7'd611 && y == 7'd434) ||
		(x == 7'd77 && y == 467) || (x == 7'd591 && y == 7'd623) || (x == 7'd601 && y == 7'd428) ||
		(x == 7'd468 && y == 7'd373) || (x == 7'd165 && y == 7'd295) || (x == 572 && y == 7'd421) ||
		(x == 7'd523 && y == 171) || (x == 7'd593 && y == 230) || (x == 7'd295 && y == 7'd596) ||
		(x == 522 && y == 7'd230) || (x == 102 && y == 7'd514) || (x == 265 && y == 477) ||
		(x == 7'd120 && y == 7'd206) || (x == 42 && y == 98) || (x == 7'd585 && y == 41) ||
		(x == 7'd317 && y == 7'd321) || (x == 7'd635 && y == 7'd412) || (x == 477 && y == 7'd97) ||
		(x == 334 && y == 7'd175) || (x == 7'd322 && y == 184) || (x == 7'd0 && y == 309) ||
		(x == 7'd615 && y == 7'd376) || (x == 243 && y == 166) || (x == 7'd2 && y == 445) ||
		(x == 398 && y == 410) || (x == 7'd274 && y == 7'd407) || (x == 342 && y == 7'd337) ||
		(x == 7'd451 && y == 571) || (x == 396 && y == 7'd270) || (x == 635 && y == 635) ||
		(x == 7'd349 && y == 207) || (x == 7'd65 && y == 247) || (x == 7'd364 && y == 7'd346) ||
		(x == 217 && y == 7'd225) || (x == 238 && y == 7'd516) || (x == 7'd192 && y == 7'd72) ||
		(x == 253 && y == 7'd181) || (x == 7'd509 && y == 7'd280) || (x == 196 && y == 7'd352) ||
		(x == 7'd308 && y == 541) || (x == 192 && y == 357) || (x == 7'd124 && y == 7'd167) ||
		(x == 140 && y == 333) || (x == 7'd31 && y == 451) || (x == 7'd282 && y == 7'd482) ||
		(x == 7'd552 && y == 444) || (x == 153 && y == 278) || (x == 7'd134 && y == 7'd516) ||
		(x == 7'd520 && y == 7'd629) || (x == 7'd432 && y == 7'd638) || (x == 303 && y == 306) ||
		(x == 7'd638 && y == 7'd334) || (x == 7'd1 && y == 143) || (x == 400 && y == 7'd613) ||
		(x == 627 && y == 314) || (x == 256 && y == 7'd508) || (x == 7'd492 && y == 7'd155) ||
		(x == 17 && y == 7'd513) || (x == 7'd588 && y == 7'd286) || (x == 7'd498 && y == 7'd423) ||
		(x == 7'd144 && y == 14) || (x == 7'd221 && y == 637) || (x == 7'd121 && y == 7'd446) ||
		(x == 214 && y == 7'd483) || (x == 44 && y == 7'd235) || (x == 306 && y == 7'd612) ||
		(x == 7'd229 && y == 7'd239) || (x == 344 && y == 7'd631) || (x == 483 && y == 7'd287) ||
		(x == 442 && y == 600) || (x == 92 && y == 7'd292) || (x == 34 && y == 7'd442) ||
		(x == 286 && y == 7'd303) || (x == 7'd402 && y == 7'd630) || (x == 7'd625 && y == 7'd449) ||
		(x == 563 && y == 7'd541) || (x == 7'd573 && y == 435) || (x == 7'd436 && y == 7'd229) ||
		(x == 240 && y == 7'd44) || (x == 7'd244 && y == 436) || (x == 7'd319 && y == 7'd141) ||
		(x == 594 && y == 7'd436) || (x == 7'd240 && y == 7'd134) || (x == 576 && y == 7'd210) ||
		(x == 7'd375 && y == 345) || (x == 7'd67 && y == 91) || (x == 7'd194 && y == 7'd167) ||
		(x == 599 && y == 599) || (x == 7'd290 && y == 640) || (x == 7'd570 && y == 626) ||
		(x == 7'd199 && y == 602) || (x == 574 && y == 409) || (x == 350 && y == 7'd409) ||
		(x == 7'd112 && y == 147) || (x == 378 && y == 386) || (x == 7'd429 && y == 7'd491) ||
		(x == 7'd289 && y == 7'd195) || (x == 7'd444 && y == 85) || (x == 7'd213 && y == 7'd260) ||
		(x == 7'd343 && y == 7'd590) || (x == 613 && y == 7'd106) || (x == 7'd343 && y == 537) ||
		(x == 7'd425 && y == 465) || (x == 7'd389 && y == 7'd203) || (x == 582 && y == 595) ||
		(x == 7'd234 && y == 405) || (x == 7'd130 && y == 7'd559) || (x == 7'd158 && y == 7'd378) ||
		(x == 7'd71 && y == 615) || (x == 7'd448 && y == 7'd93) || (x == 163 && y == 7'd212) ||
		(x == 7'd545 && y == 7'd347) || (x == 7'd54 && y == 7'd239) || (x == 7'd473 && y == 408) ||
		(x == 225 && y == 613) || (x == 508 && y == 520) || (x == 7'd489 && y == 7'd305) ||
		(x == 7'd506 && y == 7'd252) || (x == 544 && y == 369) || (x == 7'd230 && y == 298) ||
		(x == 7'd231 && y == 7'd258) || (x == 396 && y == 7'd384) || (x == 7'd259 && y == 470) ||
		(x == 276 && y == 7'd408) || (x == 7'd421 && y == 0) || (x == 7'd368 && y == 7'd27) ||
		(x == 548 && y == 410) || (x == 7'd332 && y == 306) || (x == 7'd568 && y == 7'd368) ||
		(x == 7'd176 && y == 7'd268) || (x == 7'd158 && y == 7'd429) || (x == 369 && y == 584) ||
		(x == 628 && y == 7'd74) || (x == 7'd543 && y == 7'd292) || (x == 64 && y == 7'd105) ||
		(x == 7'd468 && y == 619) || (x == 361 && y == 218) || (x == 7'd562 && y == 7'd102) ||
		(x == 233 && y == 7'd142) || (x == 7'd151 && y == 402) || (x == 151 && y == 306) ||
		(x == 7'd329 && y == 7'd144) || (x == 7'd424 && y == 7'd248) || (x == 419 && y == 386) ||
		(x == 7'd232 && y == 7'd458) || (x == 433 && y == 190) || (x == 7'd298 && y == 236) ||
		(x == 571 && y == 7'd450) || (x == 479 && y == 7'd606) || (x == 11 && y == 7'd573) ||
		(x == 384 && y == 638) || (x == 7'd394 && y == 7'd145) || (x == 7'd84 && y == 7'd248) ||
		(x == 7'd395 && y == 7'd129) || (x == 470 && y == 7'd94) || (x == 7'd89 && y == 7'd244) ||
		(x == 7'd109 && y == 7'd3) || (x == 176 && y == 310) || (x == 7'd6 && y == 7'd290) ||
		(x == 7'd426 && y == 7'd240) || (x == 345 && y == 587) || (x == 235 && y == 7'd326) ||
		(x == 361 && y == 7'd629) || (x == 7'd399 && y == 618) || (x == 7'd356 && y == 191) ||
		(x == 28 && y == 7'd390) || (x == 7'd245 && y == 186) || (x == 7'd115 && y == 385) ||
		(x == 349 && y == 282) || (x == 7'd333 && y == 7'd558) || (x == 200 && y == 7'd138) ||
		(x == 7'd580 && y == 7'd179) || (x == 7'd265 && y == 91) || (x == 189 && y == 7'd524) ||
		(x == 7'd236 && y == 334) || (x == 7'd238 && y == 201) || (x == 26 && y == 7'd310) ||
		(x == 424 && y == 7'd204) || (x == 321 && y == 7'd212) || (x == 327 && y == 7'd178) ||
		(x == 7'd206 && y == 602) || (x == 7'd340 && y == 391) || (x == 7'd138 && y == 7'd91) ||
		(x == 293 && y == 610) || (x == 7'd446 && y == 7'd248) || (x == 188 && y == 7'd29) ||
		(x == 7'd614 && y == 462) || (x == 7'd313 && y == 7'd257) || (x == 190 && y == 7'd26) ||
		(x == 312 && y == 7'd505) || (x == 7'd204 && y == 614) || (x == 7'd67 && y == 7'd524) ||
		(x == 7'd518 && y == 7'd456) || (x == 541 && y == 7'd16) || (x == 7'd184 && y == 84) ||
		(x == 7'd509 && y == 7'd195) || (x == 7'd299 && y == 7'd95) || (x == 7'd451 && y == 73) ||
		(x == 7'd275 && y == 83) || (x == 419 && y == 451) || (x == 621 && y == 622) ||
		(x == 7'd464 && y == 7'd345) || (x == 7'd491 && y == 7'd353) || (x == 7'd468 && y == 7'd372) ||
		(x == 7'd163 && y == 584) || (x == 397 && y == 598) || (x == 7'd66 && y == 7'd69) ||
		(x == 7'd499 && y == 7'd271) || (x == 313 && y == 617) || (x == 7'd220 && y == 7'd163) ||
		(x == 584 && y == 534) || (x == 267 && y == 177) || (x == 7'd400 && y == 359) ||
		(x == 167 && y == 278) || (x == 283 && y == 7'd640) || (x == 7'd450 && y == 7'd454) ||
		(x == 7'd318 && y == 7'd601) || (x == 395 && y == 7'd373) || (x == 536 && y == 7'd178) ||
		(x == 149 && y == 7'd38) || (x == 7'd210 && y == 7'd432) || (x == 7'd231 && y == 46) ||
		(x == 7'd327 && y == 7'd334) || (x == 278 && y == 7'd414) || (x == 7'd443 && y == 7'd133) ||
		(x == 7'd228 && y == 7'd621) || (x == 7'd27 && y == 7'd45) || (x == 7'd19 && y == 7'd172) ||
		(x == 7'd578 && y == 7'd632) || (x == 149 && y == 7'd78) || (x == 7'd237 && y == 237) ||
		(x == 103 && y == 7'd610) || (x == 7'd112 && y == 464) || (x == 433 && y == 477) ||
		(x == 7'd624 && y == 415) || (x == 321 && y == 338) || (x == 7'd54 && y == 432) ||
		(x == 7'd544 && y == 282) || (x == 530 && y == 7'd324) || (x == 7'd595 && y == 124) ||
		(x == 7'd568 && y == 7'd380) || (x == 487 && y == 7'd4) || (x == 190 && y == 181) ||
		(x == 7'd476 && y == 183) || (x == 7'd262 && y == 7'd268) || (x == 7'd162 && y == 7'd355) ||
		(x == 7'd297 && y == 7'd242) || (x == 155 && y == 7'd457) || (x == 7'd604 && y == 89) ||
		(x == 130 && y == 7'd158) || (x == 527 && y == 572) || (x == 7'd140 && y == 7'd599) ||
		(x == 7'd339 && y == 7'd175) || (x == 329 && y == 7'd303) || (x == 7'd345 && y == 498) ||
		(x == 7'd86 && y == 7'd274) || (x == 7'd140 && y == 330) || (x == 141 && y == 7'd83) ||
		(x == 147 && y == 7'd244) || (x == 7'd519 && y == 7'd347) || (x == 485 && y == 226) ||
		(x == 7'd340 && y == 559) || (x == 7'd188 && y == 429) || (x == 7'd451 && y == 7'd295) ||
		(x == 514 && y == 7'd557) || (x == 7'd398 && y == 7'd59) || (x == 7'd154 && y == 7'd177) ||
		(x == 58 && y == 7'd112) || (x == 7'd299 && y == 122) || (x == 524 && y == 285) ||
		(x == 7'd234 && y == 504) || (x == 7'd255 && y == 7'd27) || (x == 7'd273 && y == 7'd0) ||
		(x == 408 && y == 7'd174) || (x == 7'd97 && y == 287) || (x == 452 && y == 7'd221) ||
		(x == 7'd440 && y == 7'd626) || (x == 7'd258 && y == 7'd157) || (x == 93 && y == 7'd122) ||
		(x == 7'd573 && y == 7'd113) || (x == 575 && y == 573) || (x == 7'd119 && y == 7'd380) ||
		(x == 7'd120 && y == 7'd589) || (x == 7'd553 && y == 7'd594) || (x == 630 && y == 153) ||
		(x == 450 && y == 7'd234) || (x == 7'd587 && y == 596) || (x == 7'd234 && y == 7'd558) ||
		(x == 7'd155 && y == 7'd171) || (x == 7'd481 && y == 445) || (x == 7'd518 && y == 56) ||
		(x == 7'd229 && y == 403) || (x == 498 && y == 269) || (x == 242 && y == 541) ||
		(x == 7'd614 && y == 262) || (x == 7'd185 && y == 583) || (x == 7'd342 && y == 525) ||
		(x == 7'd598 && y == 7'd604) || (x == 7'd422 && y == 7'd235) || (x == 7'd211 && y == 7'd177) ||
		(x == 166 && y == 7'd394) || (x == 350 && y == 7'd415) || (x == 7'd348 && y == 521) ||
		(x == 272 && y == 586) || (x == 530 && y == 7'd377) || (x == 7'd180 && y == 7'd257) ||
		(x == 7'd273 && y == 7'd131) || (x == 7'd255 && y == 361) || (x == 7'd159 && y == 487) ||
		(x == 7'd561 && y == 395) || (x == 237 && y == 7'd303) || (x == 193 && y == 543) ||
		(x == 214 && y == 581) || (x == 7'd80 && y == 213) || (x == 7'd163 && y == 7'd344) ||
		(x == 7'd571 && y == 611) || (x == 7'd346 && y == 7'd370) || (x == 408 && y == 549) ||
		(x == 7'd244 && y == 75) || (x == 445 && y == 429) || (x == 597 && y == 560) ||
		(x == 7'd150 && y == 7'd411) || (x == 7'd518 && y == 7'd206) || (x == 7'd233 && y == 299) ||
		(x == 329 && y == 201) || (x == 7'd245 && y == 7'd366) || (x == 7'd605 && y == 318) ||
		(x == 7'd290 && y == 121) || (x == 7'd38 && y == 242) || (x == 237 && y == 7'd215) ||
		(x == 7'd185 && y == 530) || (x == 198 && y == 7'd368) || (x == 7'd350 && y == 7'd342) ||
		(x == 7'd531 && y == 7'd590) || (x == 7'd598 && y == 540) || (x == 229 && y == 7'd328) ||
		(x == 7'd132 && y == 174) || (x == 7'd351 && y == 7'd125) || (x == 182 && y == 7'd542) ||
		(x == 236 && y == 7'd126) || (x == 7'd151 && y == 126) || (x == 304 && y == 7'd16) ||
		(x == 7'd390 && y == 107) || (x == 7'd247 && y == 148) || (x == 7'd316 && y == 502) ||
		(x == 7'd303 && y == 7'd527) || (x == 7'd104 && y == 7'd85) || (x == 7'd97 && y == 288) ||
		(x == 254 && y == 518) || (x == 7'd201 && y == 556) || (x == 7'd434 && y == 177) ||
		(x == 7'd263 && y == 7'd55) || (x == 431 && y == 7'd615) || (x == 629 && y == 453) ||
		(x == 7'd428 && y == 500) || (x == 587 && y == 206) || (x == 7'd266 && y == 7'd464) ||
		(x == 229 && y == 501) || (x == 7'd276 && y == 7'd324) || (x == 7'd175 && y == 7'd158) ||
		(x == 229 && y == 535) || (x == 7'd634 && y == 7'd168) || (x == 539 && y == 7'd67) ||
		(x == 7'd132 && y == 7'd507) || (x == 579 && y == 461) || (x == 7'd366 && y == 7'd193) ||
		(x == 486 && y == 7'd420) || (x == 7'd268 && y == 7'd88) || (x == 7'd108 && y == 597) ||
		(x == 7'd389 && y == 7'd200) || (x == 7'd256 && y == 185) || (x == 496 && y == 7'd457) ||
		(x == 222 && y == 7'd15) || (x == 7'd305 && y == 7'd332) || (x == 7'd583 && y == 481) ||
		(x == 7'd493 && y == 7'd553) || (x == 7'd18 && y == 553) || (x == 7'd504 && y == 6) ||
		(x == 635 && y == 183) || (x == 574 && y == 7'd83) || (x == 246 && y == 7'd281) ||
		(x == 381 && y == 7'd587) || (x == 7'd520 && y == 621) || (x == 246 && y == 204) ||
		(x == 7'd620 && y == 450) || (x == 7'd470 && y == 7'd228) || (x == 428 && y == 7'd65) ||
		(x == 7'd289 && y == 449) || (x == 7'd308 && y == 7'd309) || (x == 280 && y == 7'd520) ||
		(x == 210 && y == 245) || (x == 160 && y == 7'd316) || (x == 287 && y == 429) ||
		(x == 7'd370 && y == 7'd495) || (x == 7'd41 && y == 7'd175) || (x == 7'd382 && y == 7'd130) ||
		(x == 104 && y == 7'd256) || (x == 419 && y == 354) || (x == 556 && y == 7'd208) ||
		(x == 7'd315 && y == 117) || (x == 482 && y == 7'd171) || (x == 314 && y == 268) ||
		(x == 364 && y == 335) || (x == 77 && y == 111) || (x == 7'd119 && y == 7'd521) ||
		(x == 7'd407 && y == 356) || (x == 450 && y == 7'd341) || (x == 7'd578 && y == 624) ||
		(x == 226 && y == 7'd432) || (x == 164 && y == 7'd630) || (x == 7'd273 && y == 7'd174) ||
		(x == 7'd336 && y == 7'd607) || (x == 7'd198 && y == 7'd382) || (x == 462 && y == 463) ||
		(x == 7'd136 && y == 534) || (x == 572 && y == 7'd368) || (x == 319 && y == 7'd390) ||
		(x == 298 && y == 408) || (x == 418 && y == 168) || (x == 7'd233 && y == 7'd211) ||
		(x == 363 && y == 261) || (x == 522 && y == 395) || (x == 606 && y == 7'd112) ||
		(x == 505 && y == 7'd494) || (x == 7'd322 && y == 242) || (x == 7'd239 && y == 7'd6) ||
		(x == 7'd574 && y == 7'd174) || (x == 7'd630 && y == 274) || (x == 7'd190 && y == 7'd352) ||
		(x == 7'd218 && y == 37) || (x == 7'd368 && y == 92) || (x == 26 && y == 7'd228) ||
		(x == 7'd397 && y == 173) || (x == 7'd119 && y == 494) || (x == 156 && y == 7'd598) ||
		(x == 7'd392 && y == 639) || (x == 7'd495 && y == 464) || (x == 591 && y == 350) ||
		(x == 616 && y == 293) || (x == 597 && y == 598) || (x == 7'd21 && y == 7'd381) ||
		(x == 7'd578 && y == 134) || (x == 7'd355 && y == 7'd168) || (x == 7'd584 && y == 7'd514) ||
		(x == 349 && y == 436) || (x == 444 && y == 7'd274) || (x == 606 && y == 7'd149) ||
		(x == 261 && y == 502) || (x == 269 && y == 322) || (x == 7'd501 && y == 636) ||
		(x == 207 && y == 7'd630) || (x == 7'd469 && y == 7'd248) || (x == 605 && y == 262) ||
		(x == 402 && y == 7'd85) || (x == 430 && y == 7'd248) || (x == 447 && y == 324) ||
		(x == 156 && y == 7'd562) || (x == 146 && y == 584) || (x == 7'd138 && y == 486) ||
		(x == 7'd605 && y == 7'd522) || (x == 7'd74 && y == 306) || (x == 7'd188 && y == 95) ||
		(x == 7'd78 && y == 263) || (x == 7'd322 && y == 7'd518) || (x == 7'd629 && y == 7'd609) ||
		(x == 7'd481 && y == 7'd138) || (x == 186 && y == 203) || (x == 600 && y == 7'd375) ||
		(x == 7'd485 && y == 613) || (x == 592 && y == 7'd91) || (x == 259 && y == 7'd379) ||
		(x == 443 && y == 205) || (x == 7'd356 && y == 7'd135) || (x == 7'd203 && y == 85) ||
		(x == 7'd263 && y == 328) || (x == 7'd575 && y == 7'd361) || (x == 7'd542 && y == 137) ||
		(x == 231 && y == 366) || (x == 136 && y == 7'd299) || (x == 431 && y == 577) ||
		(x == 7'd247 && y == 7'd72) || (x == 7'd222 && y == 7'd271) || (x == 7'd377 && y == 522) ||
		(x == 404 && y == 7'd378) || (x == 474 && y == 7'd507) || (x == 7'd454 && y == 7'd552) ||
		(x == 378 && y == 7'd508) || (x == 7'd122 && y == 7'd396) || (x == 281 && y == 7'd222) ||
		(x == 527 && y == 7'd68) || (x == 7'd457 && y == 17) || (x == 7'd406 && y == 7'd438) ||
		(x == 7'd448 && y == 7'd210) || (x == 7'd506 && y == 514) || (x == 281 && y == 7'd426) ||
		(x == 528 && y == 7'd394) || (x == 480 && y == 7'd13) || (x == 7'd47 && y == 123) ||
		(x == 218 && y == 268) || (x == 7'd625 && y == 7'd451) || (x == 207 && y == 7'd536) ||
		(x == 7'd633 && y == 210) || (x == 38 && y == 7'd528) || (x == 457 && y == 318) ||
		(x == 7'd130 && y == 398) || (x == 7'd233 && y == 610) || (x == 7'd499 && y == 7'd266) ||
		(x == 573 && y == 199) || (x == 553 && y == 415) || (x == 7'd20 && y == 109) ||
		(x == 326 && y == 7'd248) || (x == 628 && y == 7'd298) || (x == 7'd540 && y == 7'd423) ||
		(x == 470 && y == 451) || (x == 7'd397 && y == 501) || (x == 319 && y == 7'd631) ||
		(x == 7'd452 && y == 7'd187) || (x == 195 && y == 7'd278) || (x == 7'd88 && y == 543) ||
		(x == 188 && y == 357) || (x == 77 && y == 52) || (x == 7'd190 && y == 597) ||
		(x == 149 && y == 341) || (x == 7'd383 && y == 7'd197) || (x == 7'd412 && y == 7'd250) ||
		(x == 20 && y == 7'd266) || (x == 7'd376 && y == 7'd422) || (x == 7'd117 && y == 7'd140) ||
		(x == 597 && y == 7'd609) || (x == 630 && y == 7'd619) || (x == 527 && y == 299) ||
		(x == 597 && y == 376) || (x == 319 && y == 384) || (x == 7'd319 && y == 7'd198) ||
		(x == 7'd592 && y == 7'd327) || (x == 541 && y == 597) || (x == 7'd404 && y == 49) ||
		(x == 7'd510 && y == 7'd577) || (x == 7'd550 && y == 7'd623) || (x == 7'd41 && y == 7'd486) ||
		(x == 359 && y == 241) || (x == 7'd572 && y == 416) || (x == 314 && y == 7'd325) ||
		(x == 7'd269 && y == 7'd446) || (x == 7'd471 && y == 7'd294) || (x == 7'd184 && y == 7'd635) ||
		(x == 497 && y == 527) || (x == 203 && y == 7'd632) || (x == 7'd451 && y == 231) ||
		(x == 7'd100 && y == 559) || (x == 7'd492 && y == 412) || (x == 131 && y == 545) ||
		(x == 513 && y == 208) || (x == 7'd266 && y == 7'd622) || (x == 429 && y == 613) ||
		(x == 523 && y == 7'd20) || (x == 7'd540 && y == 7'd389) || (x == 7'd131 && y == 7'd480) ||
		(x == 279 && y == 7'd262) || (x == 7'd326 && y == 296) || (x == 7'd443 && y == 7'd239) ||
		(x == 7'd117 && y == 438) || (x == 617 && y == 7'd416) || (x == 7'd210 && y == 189) ||
		(x == 7'd41 && y == 264) || (x == 7'd187 && y == 64) || (x == 250 && y == 285) ||
		(x == 7'd485 && y == 7'd455) || (x == 7'd224 && y == 7'd465) || (x == 7'd473 && y == 7'd459) ||
		(x == 261 && y == 557) || (x == 7'd436 && y == 479) || (x == 7'd330 && y == 230) ||
		(x == 483 && y == 314) || (x == 7'd379 && y == 569) || (x == 629 && y == 272) ||
		(x == 496 && y == 7'd278) || (x == 7'd576 && y == 7'd556) || (x == 7'd228 && y == 7'd388) ||
		(x == 7'd172 && y == 623) || (x == 7'd259 && y == 7'd614) || (x == 38 && y == 7'd134) ||
		(x == 444 && y == 276) || (x == 516 && y == 549) || (x == 7'd45 && y == 62) ||
		(x == 185 && y == 552) || (x == 7'd376 && y == 7'd272) || (x == 470 && y == 7'd185) ||
		(x == 7'd589 && y == 48) || (x == 7'd245 && y == 7'd84) || (x == 7'd509 && y == 442) ||
		(x == 7'd581 && y == 7'd562) || (x == 368 && y == 532) || (x == 184 && y == 7'd120) ||
		(x == 7'd161 && y == 101) || (x == 7'd593 && y == 7'd229) || (x == 7'd565 && y == 417) ||
		(x == 7'd579 && y == 351) || (x == 179 && y == 7'd260) || (x == 7'd482 && y == 7'd403) ||
		(x == 350 && y == 7'd438) || (x == 7'd23 && y == 7'd137) || (x == 194 && y == 7'd300) ||
		(x == 421 && y == 351) || (x == 240 && y == 7'd180) || (x == 7'd41 && y == 367) ||
		(x == 424 && y == 7'd282) || (x == 7'd569 && y == 7'd584) || (x == 14 && y == 1) ||
		(x == 276 && y == 7'd625) || (x == 7'd187 && y == 617) || (x == 120 && y == 7'd215) ||
		(x == 351 && y == 7'd430) || (x == 7'd111 && y == 7'd436) || (x == 334 && y == 7'd328) ||
		(x == 7'd473 && y == 7'd134) || (x == 17 && y == 7'd291) || (x == 7'd612 && y == 299) ||
		(x == 7'd393 && y == 7'd460) || (x == 7'd59 && y == 514) || (x == 519 && y == 7'd130) ||
		(x == 7'd217 && y == 7'd208) || (x == 7'd124 && y == 7'd256) || (x == 525 && y == 7'd133) ||
		(x == 7'd378 && y == 7'd391) || (x == 432 && y == 7'd249) || (x == 7'd294 && y == 332) ||
		(x == 7'd541 && y == 236) || (x == 611 && y == 7'd533) || (x == 7'd461 && y == 7'd510) ||
		(x == 7'd72 && y == 39) || (x == 7'd135 && y == 7'd221) || (x == 7'd538 && y == 248) ||
		(x == 7'd61 && y == 547) || (x == 7'd1 && y == 146) || (x == 7'd457 && y == 7'd435) ||
		(x == 7'd492 && y == 7'd157) || (x == 7'd568 && y == 7'd196) || (x == 610 && y == 295) ||
		(x == 7'd344 && y == 507) || (x == 7'd108 && y == 7'd298) || (x == 429 && y == 7'd324) ||
		(x == 438 && y == 7'd228) || (x == 363 && y == 256) || (x == 583 && y == 162) ||
		(x == 594 && y == 561) || (x == 448 && y == 7'd276) || (x == 422 && y == 7'd390) ||
		(x == 7'd211 && y == 7'd560) || (x == 7'd140 && y == 7'd627) || (x == 7'd13 && y == 174) ||
		(x == 571 && y == 356) || (x == 178 && y == 7'd191) || (x == 7'd511 && y == 7'd406) ||
		(x == 7'd417 && y == 528) || (x == 571 && y == 7'd386) || (x == 7'd470 && y == 141) ||
		(x == 7'd581 && y == 7'd463) || (x == 380 && y == 7'd526) || (x == 7'd509 && y == 7'd277) ||
		(x == 7'd414 && y == 7'd619) || (x == 72 && y == 7'd619) || (x == 574 && y == 7'd399) ||
		(x == 7'd89 && y == 528) || (x == 7'd219 && y == 259) || (x == 7'd24 && y == 616) ||
		(x == 7'd493 && y == 282) || (x == 346 && y == 7'd507) || (x == 552 && y == 7'd134) ||
		(x == 431 && y == 7'd182) || (x == 7'd275 && y == 7'd524) || (x == 7'd121 && y == 416) ||
		(x == 492 && y == 7'd198) || (x == 7'd190 && y == 28) || (x == 7'd638 && y == 7'd171) ||
		(x == 7'd128 && y == 289) || (x == 449 && y == 283) || (x == 7'd452 && y == 618) ||
		(x == 273 && y == 7'd477) || (x == 7'd618 && y == 480) || (x == 7'd232 && y == 7'd428) ||
		(x == 7'd172 && y == 124) || (x == 272 && y == 501) || (x == 7'd56 && y == 399) ||
		(x == 7'd214 && y == 185) || (x == 7'd336 && y == 450) || (x == 7'd215 && y == 7'd17) ||
		(x == 547 && y == 290) || (x == 7'd156 && y == 447) || (x == 481 && y == 178) ||
		(x == 157 && y == 7'd185) || (x == 401 && y == 191) || (x == 7'd633 && y == 7'd233) ||
		(x == 7'd281 && y == 129) || (x == 7'd34 && y == 493) || (x == 7'd546 && y == 7'd65) ||
		(x == 593 && y == 7'd301) || (x == 7'd518 && y == 344) || (x == 492 && y == 368) ||
		(x == 7'd56 && y == 7'd573) || (x == 562 && y == 7'd174) || (x == 552 && y == 504) ||
		(x == 160 && y == 247) || (x == 7'd244 && y == 348) || (x == 7'd222 && y == 180) ||
		(x == 541 && y == 319) || (x == 7'd160 && y == 537) || (x == 7'd533 && y == 7'd264) ||
		(x == 7'd495 && y == 489) || (x == 7'd194 && y == 7'd337) || (x == 202 && y == 238) ||
		(x == 7'd255 && y == 7'd504) || (x == 7'd144 && y == 7'd599) || (x == 441 && y == 7'd293) ||
		(x == 509 && y == 7'd119) || (x == 7'd601 && y == 396) || (x == 7'd244 && y == 7'd378) ||
		(x == 422 && y == 565) || (x == 452 && y == 7'd49) || (x == 246 && y == 636) ||
		(x == 7'd484 && y == 355) || (x == 163 && y == 588) || (x == 495 && y == 7'd392) ||
		(x == 7'd405 && y == 7'd10) || (x == 264 && y == 245) || (x == 78 && y == 7'd622) ||
		(x == 452 && y == 356) || (x == 7'd431 && y == 482) || (x == 7'd194 && y == 136) ||
		(x == 465 && y == 7'd17) || (x == 7'd80 && y == 182) || (x == 7'd273 && y == 7'd260) ||
		(x == 102 && y == 7'd257) || (x == 398 && y == 561) || (x == 7'd415 && y == 229) ||
		(x == 290 && y == 560) || (x == 451 && y == 560) || (x == 635 && y == 621) ||
		(x == 7'd548 && y == 7'd388) || (x == 148 && y == 7'd145) || (x == 566 && y == 7'd493) ||
		(x == 7'd359 && y == 7'd154) || (x == 368 && y == 278) || (x == 449 && y == 446) ||
		(x == 7'd229 && y == 7'd621) || (x == 7'd175 && y == 7'd382) || (x == 519 && y == 7'd511) ||
		(x == 7'd362 && y == 7'd534) || (x == 7'd118 && y == 597) || (x == 460 && y == 149) ||
		(x == 7'd164 && y == 7'd398) || (x == 586 && y == 7'd365) || (x == 7'd376 && y == 7'd64) ||
		(x == 7'd425 && y == 13) || (x == 7'd181 && y == 7'd536) || (x == 243 && y == 7'd83) ||
		(x == 7'd447 && y == 142) || (x == 7'd388 && y == 7'd509) || (x == 7'd132 && y == 7'd543) ||
		(x == 7'd236 && y == 7'd406) || (x == 572 && y == 351) || (x == 359 && y == 7'd606) ||
		(x == 7'd294 && y == 7'd524) || (x == 7'd111 && y == 7'd65) || (x == 448 && y == 496) ||
		(x == 450 && y == 7'd229) || (x == 7'd370 && y == 7'd441) || (x == 7'd325 && y == 7'd113) ||
		(x == 7'd492 && y == 7'd25) || (x == 457 && y == 7'd42) || (x == 636 && y == 7'd573) ||
		(x == 7'd395 && y == 7'd145) || (x == 561 && y == 7'd101) || (x == 26 && y == 7'd105) ||
		(x == 7'd178 && y == 518) || (x == 7'd236 && y == 7'd248) || (x == 559 && y == 291) ||
		(x == 488 && y == 7'd314) || (x == 7'd441 && y == 164) || (x == 7'd626 && y == 7'd517) ||
		(x == 382 && y == 143) || (x == 7'd45 && y == 7'd223) || (x == 7'd292 && y == 7'd20) ||
		(x == 7'd124 && y == 7'd130) || (x == 619 && y == 331) || (x == 7'd491 && y == 86) ||
		(x == 7'd491 && y == 98) || (x == 7'd231 && y == 7'd133) || (x == 7'd375 && y == 7'd494) ||
		(x == 296 && y == 206) || (x == 7'd13 && y == 7'd570) || (x == 7'd612 && y == 289) ||
		(x == 450 && y == 144) || (x == 493 && y == 272) || (x == 615 && y == 7'd320) ||
		(x == 7'd484 && y == 603) || (x == 7'd571 && y == 151) || (x == 263 && y == 628) ||
		(x == 198 && y == 310) || (x == 308 && y == 7'd418) || (x == 7'd166 && y == 190) ||
		(x == 414 && y == 7'd16) || (x == 191 && y == 611) || (x == 507 && y == 7'd566) ||
		(x == 7'd300 && y == 75) || (x == 7'd629 && y == 7'd473) || (x == 69 && y == 7'd310) ||
		(x == 7'd414 && y == 172) || (x == 366 && y == 7'd167) || (x == 7'd514 && y == 430) ||
		(x == 7'd193 && y == 13) || (x == 7'd518 && y == 7'd360) || (x == 7'd65 && y == 7'd395) ||
		(x == 7'd553 && y == 7'd505) || (x == 7'd283 && y == 7'd617) || (x == 110 && y == 7'd156) ||
		(x == 7'd493 && y == 402) || (x == 7'd539 && y == 7'd506) || (x == 7'd273 && y == 7'd619) ||
		(x == 108 && y == 7'd427) || (x == 7'd358 && y == 7'd336) || (x == 7'd31 && y == 7'd469) ||
		(x == 7'd307 && y == 7'd132) || (x == 274 && y == 7'd383) || (x == 7'd446 && y == 67) ||
		(x == 7'd137 && y == 7'd450) || (x == 569 && y == 188) || (x == 593 && y == 7'd412) ||
		(x == 7'd131 && y == 7'd307) || (x == 208 && y == 7'd233) || (x == 7'd281 && y == 7'd363) ||
		(x == 494 && y == 7'd234) || (x == 329 && y == 316) || (x == 7'd184 && y == 465) ||
		(x == 7'd172 && y == 268) || (x == 7'd446 && y == 251) || (x == 447 && y == 212) ||
		(x == 343 && y == 254) || (x == 318 && y == 138) || (x == 413 && y == 461) ||
		(x == 7'd613 && y == 480) || (x == 433 && y == 7'd244) || (x == 21 && y == 24) ||
		(x == 259 && y == 621) || (x == 406 && y == 330) || (x == 7'd474 && y == 7'd557) ||
		(x == 7'd244 && y == 54) || (x == 627 && y == 7'd280) || (x == 7'd261 && y == 574) ||
		(x == 600 && y == 7'd192) || (x == 202 && y == 244) || (x == 7'd345 && y == 605) ||
		(x == 37 && y == 7'd500) || (x == 7'd136 && y == 7'd504) || (x == 7'd73 && y == 548) ||
		(x == 635 && y == 7'd622) || (x == 349 && y == 7'd280) || (x == 248 && y == 622) ||
		(x == 163 && y == 7'd371) || (x == 517 && y == 142) || (x == 216 && y == 7'd526) ||
		(x == 7'd263 && y == 7'd429) || (x == 7'd393 && y == 7'd235) || (x == 161 && y == 7'd481) ||
		(x == 7'd596 && y == 7'd206) || (x == 527 && y == 7'd555) || (x == 7'd110 && y == 549) ||
		(x == 257 && y == 7'd156) || (x == 7'd325 && y == 101) || (x == 230 && y == 7'd138) ||
		(x == 7'd430 && y == 7'd637) || (x == 7'd296 && y == 7'd239) || (x == 497 && y == 7'd584) ||
		(x == 7'd266 && y == 7'd335) || (x == 394 && y == 7'd185) || (x == 264 && y == 355) ||
		(x == 556 && y == 385) || (x == 253 && y == 291) || (x == 506 && y == 592) ||
		(x == 7'd392 && y == 233) || (x == 7'd253 && y == 7'd209) || (x == 7'd214 && y == 7'd172) ||
		(x == 400 && y == 7'd208) || (x == 7'd203 && y == 424) || (x == 275 && y == 495) ||
		(x == 251 && y == 7'd114) || (x == 7'd319 && y == 142) || (x == 335 && y == 414) ||
		(x == 7'd84 && y == 7'd369) || (x == 7'd177 && y == 291) || (x == 7'd454 && y == 7'd76) ||
		(x == 7'd375 && y == 7'd542) || (x == 613 && y == 7'd591) || (x == 525 && y == 368) ||
		(x == 7'd291 && y == 118) || (x == 7'd23 && y == 421) || (x == 7'd246 && y == 14) ||
		(x == 7'd96 && y == 7'd546) || (x == 467 && y == 517) || (x == 7'd224 && y == 7'd295) ||
		(x == 7'd268 && y == 621) || (x == 425 && y == 140) || (x == 7'd63 && y == 7'd501) ||
		(x == 7'd600 && y == 7'd432) || (x == 368 && y == 7'd83) || (x == 484 && y == 7'd382) ||
		(x == 7'd547 && y == 7'd212) || (x == 261 && y == 7'd472) || (x == 7'd519 && y == 7'd220) ||
		(x == 7'd465 && y == 420) || (x == 7'd488 && y == 7'd466) || (x == 7'd579 && y == 548) ||
		(x == 7'd55 && y == 7'd635) || (x == 325 && y == 7'd588) || (x == 528 && y == 7'd194) ||
		(x == 7'd637 && y == 604) || (x == 7'd193 && y == 7'd116) || (x == 7'd441 && y == 7'd251) ||
		(x == 7'd567 && y == 7'd240) || (x == 7'd638 && y == 561) || (x == 226 && y == 7'd389) ||
		(x == 295 && y == 153) || (x == 7'd339 && y == 529) || (x == 156 && y == 534) ||
		(x == 327 && y == 153) || (x == 148 && y == 7'd89) || (x == 7'd96 && y == 483) ||
		(x == 7'd446 && y == 7'd299) || (x == 7'd261 && y == 583) || (x == 229 && y == 176) ||
		(x == 324 && y == 501) || (x == 7'd203 && y == 7'd603) || (x == 7'd107 && y == 417) ||
		(x == 286 && y == 399) || (x == 417 && y == 7'd224) || (x == 498 && y == 220) ||
		(x == 345 && y == 7'd503) || (x == 7'd637 && y == 7'd538) || (x == 7'd538 && y == 51) ||
		(x == 578 && y == 368) || (x == 7'd378 && y == 436) || (x == 220 && y == 399) ||
		(x == 7'd413 && y == 7'd504) || (x == 212 && y == 7'd513) || (x == 138 && y == 7'd203) ||
		(x == 7'd432 && y == 24) || (x == 7'd273 && y == 7'd186) || (x == 7'd136 && y == 7'd182) ||
		(x == 7'd218 && y == 7'd396) || (x == 632 && y == 7'd78) || (x == 388 && y == 309) ||
		(x == 392 && y == 189) || (x == 7'd459 && y == 345) || (x == 7'd14 && y == 7'd271) ||
		(x == 7'd621 && y == 7'd473) || (x == 7'd20 && y == 362) || (x == 518 && y == 7'd230) ||
		(x == 314 && y == 7'd250) || (x == 585 && y == 347) || (x == 7'd132 && y == 7'd227) ||
		(x == 540 && y == 7'd387) || (x == 609 && y == 536) || (x == 539 && y == 7'd609) ||
		(x == 7'd135 && y == 7'd237) || (x == 7'd509 && y == 7'd374) || (x == 7'd140 && y == 7'd274) ||
		(x == 7'd414 && y == 268) || (x == 7'd286 && y == 7'd174) || (x == 7'd494 && y == 7'd323) ||
		(x == 7'd263 && y == 7'd236) || (x == 202 && y == 281) || (x == 528 && y == 7'd317) ||
		(x == 7'd398 && y == 7'd593) || (x == 296 && y == 7'd511) || (x == 508 && y == 181) ||
		(x == 7'd330 && y == 7'd178) || (x == 7'd540 && y == 564) || (x == 153 && y == 7'd563) ||
		(x == 485 && y == 227) || (x == 413 && y == 7'd115) || (x == 7'd271 && y == 7'd141) ||
		(x == 7'd566 && y == 7'd510) || (x == 7'd52 && y == 7'd479) || (x == 361 && y == 176) ||
		(x == 393 && y == 265) || (x == 552 && y == 378) || (x == 7'd627 && y == 7'd416) ||
		(x == 7'd380 && y == 593) || (x == 7'd294 && y == 7'd445) || (x == 7'd311 && y == 7'd611) ||
		(x == 7'd224 && y == 237) || (x == 7'd527 && y == 235) || (x == 7'd630 && y == 7'd472) ||
		(x == 7'd332 && y == 7'd509) || (x == 391 && y == 7'd630) || (x == 522 && y == 7'd259) ||
		(x == 7'd277 && y == 7'd580) || (x == 224 && y == 7'd186) || (x == 570 && y == 7'd467) ||
		(x == 550 && y == 264) || (x == 605 && y == 639) || (x == 7'd375 && y == 7'd519) ||
		(x == 7'd538 && y == 469) || (x == 7'd170 && y == 227) || (x == 7'd184 && y == 7'd512) ||
		(x == 7'd71 && y == 7'd40) || (x == 7'd297 && y == 7'd593) || (x == 7'd545 && y == 35) ||
		(x == 3 && y == 7'd177) || (x == 7'd603 && y == 46) || (x == 7'd418 && y == 7'd619) ||
		(x == 145 && y == 7'd139) || (x == 7'd197 && y == 7'd560) || (x == 7'd568 && y == 392) ||
		(x == 7'd246 && y == 7'd598) || (x == 7'd587 && y == 7'd305) || (x == 7'd526 && y == 7'd211) ||
		(x == 7'd282 && y == 7'd230) || (x == 262 && y == 7'd158) || (x == 7'd567 && y == 371) ||
		(x == 149 && y == 610) || (x == 153 && y == 7'd301) || (x == 7'd319 && y == 7'd142) ||
		(x == 7'd611 && y == 7'd239) || (x == 192 && y == 147) || (x == 7'd177 && y == 7'd396) ||
		(x == 7'd481 && y == 291) || (x == 464 && y == 437) || (x == 92 && y == 7'd122) ||
		(x == 7'd616 && y == 494) || (x == 122 && y == 7'd230) || (x == 137 && y == 7'd194) ||
		(x == 7'd61 && y == 7'd129) || (x == 7'd364 && y == 333) || (x == 7'd139 && y == 7'd552) ||
		(x == 7'd320 && y == 59) || (x == 7'd588 && y == 154) || (x == 530 && y == 7'd179) ||
		(x == 6 && y == 7'd555) || (x == 7'd71 && y == 7'd182) || (x == 633 && y == 171) ||
		(x == 441 && y == 7'd73) || (x == 7'd224 && y == 7'd398) || (x == 542 && y == 445) ||
		(x == 7'd517 && y == 7'd389) || (x == 620 && y == 522) || (x == 7'd572 && y == 7'd289) ||
		(x == 7'd271 && y == 82) || (x == 7'd320 && y == 7'd395) || (x == 7'd522 && y == 7'd259) ||
		(x == 7'd387 && y == 439) || (x == 7'd549 && y == 7'd491) || (x == 612 && y == 187) ||
		(x == 217 && y == 7'd557) || (x == 7'd445 && y == 7) || (x == 7'd619 && y == 7'd352) ||
		(x == 7'd30 && y == 162) || (x == 7'd505 && y == 7'd614) || (x == 180 && y == 7'd34) ||
		(x == 592 && y == 7'd527) || (x == 575 && y == 7'd416) || (x == 198 && y == 454) ||
		(x == 7'd539 && y == 148) || (x == 7'd64 && y == 7'd446) || (x == 7'd229 && y == 7'd615) ||
		(x == 429 && y == 7'd460) || (x == 7'd595 && y == 7'd215) || (x == 351 && y == 532) ||
		(x == 592 && y == 7'd495) || (x == 604 && y == 7'd143) || (x == 7'd373 && y == 7'd623) ||
		(x == 299 && y == 159) || (x == 7'd154 && y == 167) || (x == 616 && y == 471) ||
		(x == 246 && y == 7'd611) || (x == 7'd366 && y == 7'd632) || (x == 76 && y == 7'd532) ||
		(x == 562 && y == 381) || (x == 7'd434 && y == 269) || (x == 176 && y == 376) ||
		(x == 450 && y == 325) || (x == 544 && y == 7'd410) || (x == 144 && y == 239) ||
		(x == 7'd506 && y == 7'd134) || (x == 596 && y == 221) || (x == 7'd562 && y == 7'd268) ||
		(x == 7'd482 && y == 247) || (x == 7'd506 && y == 7'd206) || (x == 7'd502 && y == 7'd137) ||
		(x == 7'd590 && y == 7'd177) || (x == 408 && y == 7'd338) || (x == 347 && y == 360) ||
		(x == 250 && y == 7'd268) || (x == 149 && y == 515) || (x == 7'd455 && y == 7'd201) ||
		(x == 66 && y == 83) || (x == 401 && y == 7'd148) || (x == 7'd70 && y == 7'd571) ||
		(x == 7'd254 && y == 7'd615) || (x == 356 && y == 7'd463) || (x == 515 && y == 7'd452) ||
		(x == 7'd110 && y == 7'd142) || (x == 7'd262 && y == 7'd27) || (x == 307 && y == 541) ||
		(x == 429 && y == 7'd480) || (x == 7'd325 && y == 468) || (x == 7'd89 && y == 7'd166) ||
		(x == 219 && y == 7'd225) || (x == 7'd0 && y == 316) || (x == 584 && y == 395) ||
		(x == 202 && y == 240) || (x == 613 && y == 440) || (x == 140 && y == 7'd240) ||
		(x == 7'd148 && y == 7'd547) || (x == 7'd105 && y == 308) || (x == 7'd533 && y == 7'd250) ||
		(x == 127 && y == 7'd590) || (x == 160 && y == 588) || (x == 633 && y == 433) ||
		(x == 348 && y == 7'd194) || (x == 68 && y == 7'd142) || (x == 7'd453 && y == 576) ||
		(x == 437 && y == 7'd255) || (x == 559 && y == 189) || (x == 160 && y == 559) ||
		(x == 7'd255 && y == 106) || (x == 166 && y == 616) || (x == 274 && y == 7'd125) ||
		(x == 7'd50 && y == 545) || (x == 7'd467 && y == 7'd67) || (x == 386 && y == 7'd619) ||
		(x == 634 && y == 479) || (x == 417 && y == 7'd203) || (x == 7'd125 && y == 7'd378) ||
		(x == 7'd497 && y == 7'd369) || (x == 7'd291 && y == 546) || (x == 493 && y == 7'd547) ||
		(x == 7'd371 && y == 450) || (x == 361 && y == 7'd134) || (x == 7'd540 && y == 7'd307) ||
		(x == 7'd327 && y == 286) || (x == 7'd491 && y == 368) || (x == 7'd519 && y == 185) ||
		(x == 337 && y == 517) || (x == 579 && y == 7'd526) || (x == 7'd366 && y == 251) ||
		(x == 507 && y == 7'd392) || (x == 306 && y == 7'd524) || (x == 515 && y == 7'd409) ||
		(x == 577 && y == 468) || (x == 306 && y == 557) || (x == 7'd139 && y == 7'd370) ||
		(x == 7'd552 && y == 332) || (x == 369 && y == 7'd252) || (x == 7'd511 && y == 7'd578) ||
		(x == 219 && y == 7'd186) || (x == 7'd413 && y == 7'd254) || (x == 476 && y == 7'd168) ||
		(x == 7'd165 && y == 7'd539) || (x == 7'd302 && y == 194) || (x == 7'd311 && y == 586) ||
		(x == 7'd353 && y == 7'd269) || (x == 7'd636 && y == 7'd373) || (x == 7'd184 && y == 7'd622) ||
		(x == 521 && y == 7'd93) || (x == 7'd282 && y == 145) || (x == 286 && y == 600) ||
		(x == 7'd235 && y == 7'd244) || (x == 100 && y == 7'd403) || (x == 457 && y == 7'd502) ||
		(x == 7'd545 && y == 7'd276) || (x == 7'd130 && y == 7'd518) || (x == 441 && y == 393) ||
		(x == 329 && y == 291) || (x == 638 && y == 380) || (x == 7'd544 && y == 7'd248) ||
		(x == 6 && y == 120) || (x == 7'd529 && y == 7'd249) || (x == 225 && y == 7'd278) ||
		(x == 7'd220 && y == 7'd418) || (x == 7'd6 && y == 295) || (x == 29 && y == 7'd547) ||
		(x == 7'd530 && y == 400) || (x == 505 && y == 7'd458) || (x == 294 && y == 230) ||
		(x == 7'd44 && y == 430) || (x == 599 && y == 230) || (x == 7'd366 && y == 38) ||
		(x == 7'd438 && y == 341) || (x == 7'd192 && y == 602) || (x == 561 && y == 551) ||
		(x == 7'd327 && y == 7'd80) || (x == 397 && y == 7'd504) || (x == 7'd497 && y == 7'd550) ||
		(x == 7'd451 && y == 7'd269) || (x == 7'd550 && y == 477) || (x == 535 && y == 7'd73) ||
		(x == 304 && y == 7'd585) || (x == 7'd638 && y == 7'd174) || (x == 7'd338 && y == 7'd250) ||
		(x == 560 && y == 217) || (x == 476 && y == 355) || (x == 7'd578 && y == 41) ||
		(x == 458 && y == 154) || (x == 7'd611 && y == 536) || (x == 7'd185 && y == 542) ||
		(x == 7'd113 && y == 56) || (x == 149 && y == 7'd552) || (x == 627 && y == 215) ||
		(x == 7'd379 && y == 7'd553) || (x == 252 && y == 613) || (x == 7'd332 && y == 575) ||
		(x == 290 && y == 151) || (x == 7'd161 && y == 7'd469) || (x == 216 && y == 7'd100) ||
		(x == 7'd81 && y == 404) || (x == 7'd531 && y == 7'd578) || (x == 57 && y == 7'd115) ||
		(x == 295 && y == 7'd292) || (x == 7'd86 && y == 7'd518) || (x == 7'd98 && y == 436) ||
		(x == 288 && y == 7'd278) || (x == 199 && y == 7'd369) || (x == 286 && y == 383) ||
		(x == 7'd108 && y == 145) || (x == 387 && y == 7'd323) || (x == 7'd620 && y == 7'd530) ||
		(x == 7'd563 && y == 594) || (x == 7'd270 && y == 7'd366) || (x == 599 && y == 218) ||
		(x == 7'd421 && y == 592) || (x == 541 && y == 362) || (x == 514 && y == 187) ||
		(x == 157 && y == 194) || (x == 7'd415 && y == 7'd122) || (x == 628 && y == 7'd408) ||
		(x == 7'd618 && y == 7'd384) || (x == 193 && y == 293) || (x == 129 && y == 7'd360) ||
		(x == 7'd298 && y == 7'd39) || (x == 7'd605 && y == 7'd416) || (x == 7'd424 && y == 7'd553) ||
		(x == 7'd141 && y == 234) || (x == 231 && y == 443) || (x == 7'd342 && y == 7'd355) ||
		(x == 7'd550 && y == 7'd241) || (x == 7'd455 && y == 397) || (x == 7'd380 && y == 7'd157) ||
		(x == 550 && y == 7'd410) || (x == 7'd98 && y == 7'd382) || (x == 7'd261 && y == 572) ||
		(x == 195 && y == 7'd275) || (x == 7'd523 && y == 150) || (x == 169 && y == 7'd152) ||
		(x == 267 && y == 7'd458) || (x == 7'd560 && y == 320) || (x == 7'd298 && y == 7'd465) ||
		(x == 630 && y == 431) || (x == 7'd308 && y == 7'd515) || (x == 223 && y == 7'd566) ||
		(x == 7'd298 && y == 7'd598) || (x == 7'd406 && y == 7'd453) || (x == 563 && y == 7'd27) ||
		(x == 171 && y == 392) || (x == 7'd373 && y == 562) || (x == 7'd498 && y == 7'd378) ||
		(x == 352 && y == 7'd316) || (x == 7'd96 && y == 7'd16) || (x == 500 && y == 7'd624) ||
		(x == 238 && y == 408) || (x == 7'd484 && y == 7'd264) || (x == 371 && y == 292) ||
		(x == 7'd323 && y == 276) || (x == 7'd265 && y == 118) || (x == 7'd59 && y == 7'd105) ||
		(x == 7'd607 && y == 333) || (x == 381 && y == 518) || (x == 7'd396 && y == 351) ||
		(x == 364 && y == 7'd634) || (x == 581 && y == 7'd381) || (x == 192 && y == 7'd532) ||
		(x == 620 && y == 179) || (x == 7'd614 && y == 7'd108) || (x == 7'd392 && y == 7'd516) ||
		(x == 60 && y == 7'd195) || (x == 545 && y == 7'd151) || (x == 7'd392 && y == 7'd534) ||
		(x == 185 && y == 406) || (x == 457 && y == 247) || (x == 503 && y == 421) ||
		(x == 244 && y == 7'd606) || (x == 7'd491 && y == 7'd555) || (x == 536 && y == 7'd230) ||
		(x == 7'd305 && y == 142) || (x == 7'd527 && y == 7'd109) || (x == 7'd275 && y == 7'd286) ||
		(x == 367 && y == 7'd180) || (x == 269 && y == 7'd249) || (x == 7'd466 && y == 373) ||
		(x == 583 && y == 7'd562) || (x == 119 && y == 87) || (x == 7'd211 && y == 7'd633) ||
		(x == 7'd110 && y == 183) || (x == 7'd280 && y == 7'd27) || (x == 173 && y == 283) ||
		(x == 75 && y == 126) || (x == 7'd537 && y == 7'd125) || (x == 7'd200 && y == 7'd260) ||
		(x == 482 && y == 7'd599) || (x == 7'd451 && y == 405) || (x == 7'd634 && y == 7'd411) ||
		(x == 7'd118 && y == 359) || (x == 7'd509 && y == 7'd131) || (x == 396 && y == 232) ||
		(x == 344 && y == 7'd619) || (x == 7'd576 && y == 7'd427) || (x == 7'd380 && y == 7'd483) ||
		(x == 7'd372 && y == 7'd576) || (x == 7'd457 && y == 7'd352) || (x == 230 && y == 7'd576) ||
		(x == 584 && y == 7'd447) || (x == 597 && y == 130) || (x == 3 && y == 7'd25) ||
		(x == 373 && y == 529) || (x == 277 && y == 7'd634) || (x == 7'd417 && y == 7'd184) ||
		(x == 7'd128 && y == 142) || (x == 380 && y == 390) || (x == 7'd143 && y == 7'd450) ||
		(x == 283 && y == 7'd292) || (x == 7'd34 && y == 378) || (x == 7'd110 && y == 7'd373) ||
		(x == 461 && y == 185) || (x == 218 && y == 7'd251) || (x == 7'd305 && y == 236) ||
		(x == 163 && y == 7'd528) || (x == 389 && y == 7'd30) || (x == 564 && y == 225) ||
		(x == 334 && y == 7'd626) || (x == 356 && y == 514) || (x == 7'd635 && y == 7'd298) ||
		(x == 7'd98 && y == 7'd488) || (x == 7'd34 && y == 558) || (x == 130 && y == 460) ||
		(x == 7'd294 && y == 7'd71) || (x == 624 && y == 7'd99) || (x == 7'd357 && y == 7'd532) ||
		(x == 609 && y == 7'd288) || (x == 199 && y == 7'd500) || (x == 309 && y == 7'd373) ||
		(x == 7'd254 && y == 7'd554) || (x == 522 && y == 171) || (x == 7'd353 && y == 392) ||
		(x == 143 && y == 7'd117) || (x == 589 && y == 159) || (x == 7'd451 && y == 188) ||
		(x == 7'd534 && y == 147) || (x == 7'd231 && y == 7'd556) || (x == 7'd533 && y == 7'd438) ||
		(x == 113 && y == 7'd452) || (x == 103 && y == 7'd540) || (x == 240 && y == 175) ||
		(x == 535 && y == 228) || (x == 7'd180 && y == 397) || (x == 578 && y == 7'd516) ||
		(x == 235 && y == 472) || (x == 7'd147 && y == 7'd566) || (x == 354 && y == 7'd202) ||
		(x == 7'd364 && y == 7'd384) || (x == 7'd405 && y == 7'd417) || (x == 611 && y == 7'd329) ||
		(x == 7'd508 && y == 7'd446) || (x == 7'd423 && y == 492) || (x == 216 && y == 132) ||
		(x == 7'd462 && y == 160) || (x == 7'd247 && y == 7'd141) || (x == 7'd375 && y == 7'd126) ||
		(x == 47 && y == 105) || (x == 330 && y == 363) || (x == 7'd491 && y == 7'd339) ||
		(x == 7'd200 && y == 7'd184) || (x == 7'd297 && y == 7'd538) || (x == 7'd493 && y == 7'd609) ||
		(x == 7'd600 && y == 7'd433) || (x == 7'd349 && y == 556) || (x == 534 && y == 512) ||
		(x == 144 && y == 7'd401) || (x == 139 && y == 155) || (x == 375 && y == 7'd43) ||
		(x == 222 && y == 249) || (x == 249 && y == 152) || (x == 7'd605 && y == 7'd621) ||
		(x == 7'd459 && y == 7'd617) || (x == 556 && y == 7'd174) || (x == 109 && y == 7'd474) ||
		(x == 7'd467 && y == 7'd120) || (x == 529 && y == 348) || (x == 7'd389 && y == 46) ||
		(x == 575 && y == 7'd425) || (x == 266 && y == 145) || (x == 7'd633 && y == 121) ||
		(x == 7'd240 && y == 7'd296) || (x == 7'd633 && y == 7'd231) || (x == 506 && y == 7'd45) ||
		(x == 7'd429 && y == 328) || (x == 7'd314 && y == 363) || (x == 219 && y == 7'd506) ||
		(x == 7'd533 && y == 551) || (x == 118 && y == 7'd507) || (x == 7'd354 && y == 7'd363) ||
		(x == 570 && y == 7'd129) || (x == 346 && y == 7'd448) || (x == 155 && y == 7'd297) ||
		(x == 635 && y == 7'd517) || (x == 7'd9 && y == 7'd278) || (x == 7'd490 && y == 7'd338) ||
		(x == 176 && y == 7'd289) || (x == 7'd239 && y == 7'd453) || (x == 7'd515 && y == 7'd542) ||
		(x == 7'd422 && y == 7'd141) || (x == 7'd255 && y == 7'd554) || (x == 237 && y == 543) ||
		(x == 7'd480 && y == 612) || (x == 142 && y == 7'd126) || (x == 7'd197 && y == 184) ||
		(x == 7'd366 && y == 133) || (x == 410 && y == 134) || (x == 275 && y == 7'd470) ||
		(x == 455 && y == 7'd560) || (x == 7'd314 && y == 7'd577) || (x == 241 && y == 475) ||
		(x == 7'd247 && y == 7'd608) || (x == 7'd137 && y == 7'd514) || (x == 7'd216 && y == 7'd378) ||
		(x == 7'd222 && y == 7'd507) || (x == 250 && y == 431) || (x == 179 && y == 165) ||
		(x == 7'd441 && y == 151) || (x == 521 && y == 527) || (x == 7'd490 && y == 385) ||
		(x == 7'd496 && y == 7'd562) || (x == 7'd408 && y == 7'd541) || (x == 507 && y == 201) ||
		(x == 106 && y == 7'd121) || (x == 7'd368 && y == 275) || (x == 226 && y == 215) ||
		(x == 448 && y == 7'd435) || (x == 601 && y == 442) || (x == 7'd124 && y == 7'd449) ||
		(x == 7'd637 && y == 7'd448) || (x == 7'd360 && y == 7'd242) || (x == 7'd582 && y == 7'd586) ||
		(x == 20 && y == 7'd281) || (x == 544 && y == 490) || (x == 630 && y == 7'd210) ||
		(x == 7'd243 && y == 129) || (x == 149 && y == 388) || (x == 7'd316 && y == 7'd3) ||
		(x == 376 && y == 363) || (x == 7'd324 && y == 615) || (x == 301 && y == 7'd533) ||
		(x == 185 && y == 413) || (x == 374 && y == 7'd121) || (x == 7'd535 && y == 333) ||
		(x == 7'd501 && y == 195) || (x == 306 && y == 7'd532) || (x == 7'd204 && y == 7'd610) ||
		(x == 476 && y == 7'd363) || (x == 184 && y == 7'd375) || (x == 457 && y == 487) ||
		(x == 513 && y == 7'd618) || (x == 532 && y == 517) || (x == 7'd69 && y == 576) ||
		(x == 7'd422 && y == 7'd453) || (x == 7'd247 && y == 7'd506) || (x == 602 && y == 228) ||
		(x == 7'd318 && y == 278) || (x == 7'd68 && y == 550) || (x == 7'd43 && y == 7'd119) ||
		(x == 316 && y == 516) || (x == 7'd388 && y == 628) || (x == 151 && y == 502) ||
		(x == 7'd389 && y == 7'd312) || (x == 7'd412 && y == 7'd427) || (x == 468 && y == 7'd570) ||
		(x == 7'd625 && y == 7'd131) || (x == 29 && y == 52) || (x == 98 && y == 7'd286) ||
		(x == 7'd594 && y == 140) || (x == 313 && y == 7'd435) || (x == 209 && y == 187) ||
		(x == 7'd266 && y == 7'd314) || (x == 7'd267 && y == 129) || (x == 559 && y == 7'd176) ||
		(x == 7'd293 && y == 2) || (x == 182 && y == 250) || (x == 7'd346 && y == 7'd391) ||
		(x == 104 && y == 7'd632) || (x == 639 && y == 227) || (x == 357 && y == 200) ||
		(x == 7'd579 && y == 206) || (x == 311 && y == 405) || (x == 336 && y == 443) ||
		(x == 7'd202 && y == 186) || (x == 7'd282 && y == 7'd638) || (x == 480 && y == 7'd280) ||
		(x == 7'd350 && y == 408) || (x == 285 && y == 7'd503) || (x == 167 && y == 214) ||
		(x == 7'd147 && y == 7'd503) || (x == 66 && y == 7'd163) || (x == 326 && y == 593) ||
		(x == 311 && y == 7'd30) || (x == 438 && y == 7'd346) || (x == 7'd563 && y == 296) ||
		(x == 455 && y == 7'd334) || (x == 118 && y == 7'd253) || (x == 12 && y == 7'd528) ||
		(x == 300 && y == 354) || (x == 7'd533 && y == 7'd29) || (x == 7'd527 && y == 7'd547) ||
		(x == 621 && y == 364) || (x == 7'd475 && y == 546) || (x == 7'd234 && y == 264) ||
		(x == 7'd333 && y == 7'd240) || (x == 7'd327 && y == 7'd169) || (x == 7'd618 && y == 296) ||
		(x == 487 && y == 7'd496) || (x == 7'd392 && y == 7'd409) || (x == 7'd578 && y == 365) ||
		(x == 7'd353 && y == 505) || (x == 7'd521 && y == 7'd146) || (x == 7'd465 && y == 7'd350) ||
		(x == 91 && y == 7'd253) || (x == 7'd318 && y == 455) || (x == 208 && y == 7'd321) ||
		(x == 617 && y == 7'd10) || (x == 7'd271 && y == 357) || (x == 15 && y == 7'd278) ||
		(x == 7'd624 && y == 7'd514) || (x == 7'd335 && y == 7'd512) || (x == 7'd122 && y == 7'd29) ||
		(x == 7'd112 && y == 129) || (x == 73 && y == 7'd398) || (x == 7'd193 && y == 370) ||
		(x == 239 && y == 175) || (x == 7'd189 && y == 7'd342) || (x == 468 && y == 7'd427) ||
		(x == 7'd172 && y == 7'd482) || (x == 171 && y == 7'd270) || (x == 7'd379 && y == 7'd488) ||
		(x == 7'd231 && y == 433) || (x == 189 && y == 7'd244) || (x == 382 && y == 515) ||
		(x == 7'd381 && y == 66) || (x == 604 && y == 7'd137) || (x == 7'd432 && y == 485) ||
		(x == 7'd485 && y == 108) || (x == 7'd453 && y == 7'd481) || (x == 531 && y == 7'd566) ||
		(x == 7'd190 && y == 7'd105) || (x == 562 && y == 478) || (x == 222 && y == 339) ||
		(x == 179 && y == 7'd508) || (x == 237 && y == 144) || (x == 7'd408 && y == 271) ||
		(x == 211 && y == 7'd557) || (x == 383 && y == 7'd212) || (x == 7'd15 && y == 561) ||
		(x == 420 && y == 317) || (x == 150 && y == 622) || (x == 315 && y == 7'd436) ||
		(x == 186 && y == 7'd366) || (x == 367 && y == 275) || (x == 313 && y == 7'd90) ||
		(x == 99 && y == 17) || (x == 330 && y == 141) || (x == 205 && y == 7'd34) ||
		(x == 7'd530 && y == 108) || (x == 345 && y == 356) || (x == 400 && y == 7'd424) ||
		(x == 7'd205 && y == 579) || (x == 9 && y == 7'd525) || (x == 386 && y == 492) ||
		(x == 7'd580 && y == 7'd455) || (x == 246 && y == 292) || (x == 7'd245 && y == 7'd166) ||
		(x == 7'd275 && y == 7'd451) || (x == 7'd456 && y == 7'd622) || (x == 151 && y == 444) ||
		(x == 7'd614 && y == 7'd253) || (x == 7'd198 && y == 7'd167) || (x == 7'd597 && y == 179) ||
		(x == 244 && y == 7'd140) || (x == 7'd19 && y == 480) || (x == 7'd323 && y == 7'd550) ||
		(x == 7'd420 && y == 380) || (x == 7'd95 && y == 7'd547) || (x == 7'd311 && y == 608) ||
		(x == 293 && y == 598) || (x == 616 && y == 631) || (x == 7'd288 && y == 7'd258) ||
		(x == 55 && y == 7'd489) || (x == 184 && y == 7'd89) || (x == 389 && y == 627) ||
		(x == 7'd616 && y == 7'd631) || (x == 442 && y == 7'd417) || (x == 471 && y == 410) ||
		(x == 551 && y == 7'd509) || (x == 7'd177 && y == 501) || (x == 421 && y == 576) ||
		(x == 390 && y == 311) || (x == 300 && y == 7'd308) || (x == 7'd628 && y == 7'd381) ||
		(x == 233 && y == 7'd124) || (x == 7'd165 && y == 7'd471) || (x == 7'd255 && y == 398) ||
		(x == 7'd355 && y == 510) || (x == 361 && y == 264) || (x == 7'd560 && y == 220) ||
		(x == 7'd365 && y == 7'd580) || (x == 7'd348 && y == 388) || (x == 354 && y == 391) ||
		(x == 7'd187 && y == 7'd314) || (x == 7'd554 && y == 393) || (x == 271 && y == 149) ||
		(x == 164 && y == 7'd151) || (x == 7'd556 && y == 7'd632) || (x == 173 && y == 324) ||
		(x == 148 && y == 184) || (x == 533 && y == 7'd441) || (x == 427 && y == 7'd325) ||
		(x == 584 && y == 7'd341) || (x == 7'd395 && y == 7'd219) || (x == 505 && y == 7'd636) ||
		(x == 435 && y == 7'd74) || (x == 7'd539 && y == 605) || (x == 7'd523 && y == 406) ||
		(x == 7'd269 && y == 7'd59) || (x == 7'd321 && y == 367) || (x == 7'd581 && y == 7'd516) ||
		(x == 612 && y == 279) || (x == 7'd175 && y == 7'd138) || (x == 596 && y == 7'd83) ||
		(x == 474 && y == 507) || (x == 254 && y == 7'd628) || (x == 593 && y == 192) ||
		(x == 7'd407 && y == 7'd7) || (x == 7'd525 && y == 401) || (x == 7'd616 && y == 112) ||
		(x == 7'd413 && y == 7'd303) || (x == 7'd535 && y == 335) || (x == 292 && y == 7'd23) ||
		(x == 7'd372 && y == 7'd107) || (x == 567 && y == 352) || (x == 7'd4 && y == 46) ||
		(x == 7'd126 && y == 528) || (x == 7'd465 && y == 7'd130) || (x == 155 && y == 296) ||
		(x == 7'd449 && y == 564) || (x == 609 && y == 7'd456) || (x == 399 && y == 505) ||
		(x == 7'd136 && y == 26) || (x == 7'd19 && y == 7'd287) || (x == 278 && y == 7'd300) ||
		(x == 555 && y == 491) || (x == 7'd565 && y == 7'd328) || (x == 7'd562 && y == 381) ||
		(x == 7'd501 && y == 7'd62) || (x == 7'd265 && y == 385) || (x == 10 && y == 7'd119) ||
		(x == 529 && y == 7'd322) || (x == 7'd143 && y == 7'd277) || (x == 7'd401 && y == 7'd160) ||
		(x == 201 && y == 407) || (x == 431 && y == 7'd364) || (x == 7'd106 && y == 299) ||
		(x == 392 && y == 188) || (x == 268 && y == 7'd391) || (x == 309 && y == 7'd46) ||
		(x == 7'd173 && y == 7'd524) || (x == 7'd556 && y == 7'd633) || (x == 482 && y == 7'd112) ||
		(x == 193 && y == 7'd518) || (x == 7'd148 && y == 638) || (x == 7'd581 && y == 7'd593) ||
		(x == 241 && y == 192) || (x == 7'd602 && y == 7'd306) || (x == 307 && y == 7'd13) ||
		(x == 7'd274 && y == 7'd180) || (x == 7'd347 && y == 512) || (x == 186 && y == 7'd541) ||
		(x == 7'd350 && y == 7'd270) || (x == 7'd508 && y == 7'd184) || (x == 309 && y == 7'd349) ||
		(x == 558 && y == 7'd111) || (x == 7'd100 && y == 225) || (x == 7'd408 && y == 7'd388) ||
		(x == 565 && y == 214) || (x == 472 && y == 7'd74) || (x == 430 && y == 7'd243) ||
		(x == 7'd500 && y == 555) || (x == 513 && y == 360) || (x == 7'd559 && y == 7'd331) ||
		(x == 7'd582 && y == 7'd297) || (x == 606 && y == 299) || (x == 345 && y == 7'd619) ||
		(x == 7'd494 && y == 94) || (x == 7'd0 && y == 553) || (x == 7'd355 && y == 7'd262) ||
		(x == 7'd137 && y == 7'd311) || (x == 571 && y == 153) || (x == 41 && y == 7'd420) ||
		(x == 477 && y == 7'd213) || (x == 26 && y == 7'd282) || (x == 220 && y == 551) ||
		(x == 518 && y == 587) || (x == 7'd242 && y == 347) || (x == 347 && y == 7'd193) ||
		(x == 7'd176 && y == 547) || (x == 7'd3 && y == 287) || (x == 7'd290 && y == 7'd318) ||
		(x == 7'd504 && y == 7'd416) || (x == 133 && y == 282) || (x == 7'd86 && y == 167) ||
		(x == 239 && y == 486) || (x == 7'd65 && y == 162) || (x == 271 && y == 353) ||
		(x == 7'd544 && y == 7'd634) || (x == 7'd420 && y == 7'd85) || (x == 7'd211 && y == 488) ||
		(x == 44 && y == 7'd395) || (x == 7'd446 && y == 7'd577) || (x == 106 && y == 7'd274) ||
		(x == 7'd607 && y == 7'd522) || (x == 7'd30 && y == 7'd248) || (x == 7'd143 && y == 7'd209) ||
		(x == 7'd77 && y == 598) || (x == 7'd558 && y == 445) || (x == 7'd241 && y == 7'd479) ||
		(x == 470 && y == 605) || (x == 185 && y == 410) || (x == 7'd423 && y == 379) ||
		(x == 487 && y == 177) || (x == 7'd267 && y == 348) || (x == 7'd570 && y == 7'd228) ||
		(x == 7'd125 && y == 7'd372) || (x == 7'd115 && y == 7'd197) || (x == 585 && y == 7'd426) ||
		(x == 7'd193 && y == 7'd374) || (x == 7'd380 && y == 7'd503) || (x == 247 && y == 7'd353) ||
		(x == 237 && y == 378) || (x == 316 && y == 7'd393) || (x == 7'd30 && y == 623) ||
		(x == 394 && y == 7'd154) || (x == 7'd585 && y == 38) || (x == 416 && y == 236) ||
		(x == 7'd541 && y == 7'd132) || (x == 7'd383 && y == 7'd487) || (x == 7'd596 && y == 7'd249) ||
		(x == 7'd364 && y == 419) || (x == 384 && y == 552) || (x == 7'd560 && y == 8) ||
		(x == 538 && y == 7'd60) || (x == 7'd473 && y == 482) || (x == 7'd396 && y == 7'd256) ||
		(x == 7'd101 && y == 604) || (x == 7'd351 && y == 7'd177) || (x == 427 && y == 603) ||
		(x == 7'd15 && y == 7'd183) || (x == 227 && y == 7'd141) || (x == 448 && y == 520) ||
		(x == 201 && y == 227) || (x == 7'd559 && y == 171) || (x == 7'd146 && y == 7'd197) ||
		(x == 31 && y == 7'd256) || (x == 125 && y == 7'd614) || (x == 269 && y == 184) ||
		(x == 532 && y == 201) || (x == 343 && y == 364) || (x == 7'd546 && y == 7'd469) ||
		(x == 7'd459 && y == 7'd148) || (x == 564 && y == 7'd596) || (x == 297 && y == 392) ||
		(x == 7'd511 && y == 7'd257) || (x == 7'd229 && y == 7'd170) || (x == 7'd244 && y == 213) ||
		(x == 7'd635 && y == 139) || (x == 7'd148 && y == 7'd431) || (x == 7'd209 && y == 7'd199) ||
		(x == 239 && y == 7'd618) || (x == 270 && y == 329) || (x == 7'd466 && y == 7'd309) ||
		(x == 7'd144 && y == 7'd342) || (x == 7'd627 && y == 88) || (x == 7'd451 && y == 283) ||
		(x == 7'd41 && y == 7'd629) || (x == 7'd511 && y == 7'd403) || (x == 7'd152 && y == 7'd412) ||
		(x == 288 && y == 148) || (x == 355 && y == 7'd446) || (x == 339 && y == 7'd202) ||
		(x == 7'd143 && y == 254) || (x == 385 && y == 514) || (x == 480 && y == 540) ||
		(x == 7'd581 && y == 186) || (x == 543 && y == 7'd584) || (x == 7'd377 && y == 573) ||
		(x == 7'd464 && y == 7'd470) || (x == 583 && y == 7'd139) || (x == 7'd13 && y == 164) ||
		(x == 7'd442 && y == 7'd340) || (x == 189 && y == 398) || (x == 7'd484 && y == 299) ||
		(x == 280 && y == 335) || (x == 490 && y == 477) || (x == 7'd1 && y == 502) ||
		(x == 7'd239 && y == 7'd157) || (x == 196 && y == 7'd417) || (x == 7'd600 && y == 7'd588) ||
		(x == 7'd404 && y == 7'd302) || (x == 207 && y == 7'd141) || (x == 7'd586 && y == 7'd402) ||
		(x == 7'd454 && y == 7'd209) || (x == 7'd426 && y == 7'd376) || (x == 121 && y == 7'd185) ||
		(x == 7'd407 && y == 7'd636) || (x == 634 && y == 233) || (x == 28 && y == 7'd252) ||
		(x == 367 && y == 573) || (x == 369 && y == 7'd43) || (x == 7'd501 && y == 7'd226) ||
		(x == 7'd271 && y == 7'd14) || (x == 483 && y == 7'd201) || (x == 7'd419 && y == 7'd342) ||
		(x == 596 && y == 7'd337) || (x == 7'd148 && y == 7'd377) || (x == 601 && y == 7'd241) ||
		(x == 7'd583 && y == 7'd518) || (x == 570 && y == 630) || (x == 7'd247 && y == 7'd526) ||
		(x == 423 && y == 590) || (x == 190 && y == 7'd189) || (x == 7'd601 && y == 7'd137) ||
		(x == 7'd16 && y == 36) || (x == 7'd577 && y == 7'd6) || (x == 278 && y == 7'd34) ||
		(x == 487 && y == 7'd489) || (x == 470 && y == 7'd596) || (x == 561 && y == 492) ||
		(x == 137 && y == 7'd462) || (x == 382 && y == 391) || (x == 536 && y == 431) ||
		(x == 417 && y == 7'd497) || (x == 409 && y == 7'd399) || (x == 526 && y == 458) ||
		(x == 7'd426 && y == 7'd29) || (x == 7'd574 && y == 7'd122) || (x == 7'd230 && y == 7'd468) ||
		(x == 7'd259 && y == 7'd390) || (x == 7'd160 && y == 66) || (x == 409 && y == 164) ||
		(x == 7'd544 && y == 269) || (x == 7'd517 && y == 7'd563) || (x == 7'd628 && y == 7'd390) ||
		(x == 7'd445 && y == 7'd401) || (x == 7'd229 && y == 7'd296) || (x == 272 && y == 7'd369) ||
		(x == 295 && y == 444) || (x == 7'd350 && y == 7'd112) || (x == 7'd125 && y == 7'd191) ||
		(x == 7'd27 && y == 309) || (x == 7'd268 && y == 7'd163) || (x == 164 && y == 252) ||
		(x == 292 && y == 7'd60) || (x == 7'd82 && y == 7'd197) || (x == 7'd553 && y == 311) ||
		(x == 7'd550 && y == 7'd598) || (x == 7'd600 && y == 7'd373) || (x == 7'd273 && y == 7'd240) ||
		(x == 15 && y == 7'd536) || (x == 207 && y == 392) || (x == 7'd628 && y == 421) ||
		(x == 512 && y == 7'd118) || (x == 519 && y == 7'd67) || (x == 7'd286 && y == 388) ||
		(x == 239 && y == 588) || (x == 7'd204 && y == 529) || (x == 7'd375 && y == 7'd12) ||
		(x == 370 && y == 7'd523) || (x == 7'd134 && y == 7'd449) || (x == 442 && y == 138) ||
		(x == 497 && y == 7'd414) || (x == 7'd441 && y == 7'd515) || (x == 7'd341 && y == 7'd206) ||
		(x == 160 && y == 569) || (x == 7'd374 && y == 7'd363) || (x == 124 && y == 7'd518) ||
		(x == 7'd149 && y == 569) || (x == 7'd500 && y == 7'd217) || (x == 7'd249 && y == 506) ||
		(x == 7'd294 && y == 443) || (x == 193 && y == 425) || (x == 427 && y == 7'd464) ||
		(x == 7'd595 && y == 7'd628) || (x == 7'd533 && y == 231) || (x == 599 && y == 7'd16) ||
		(x == 260 && y == 485) || (x == 7'd526 && y == 326) || (x == 7'd459 && y == 7'd271) ||
		(x == 7'd413 && y == 7'd258) || (x == 59 && y == 7'd210) || (x == 393 && y == 429) ||
		(x == 7'd260 && y == 7'd435) || (x == 7'd564 && y == 529) || (x == 7'd242 && y == 7'd520) ||
		(x == 384 && y == 326) || (x == 7'd466 && y == 7'd131) || (x == 7'd53 && y == 176) ||
		(x == 7'd27 && y == 210) || (x == 7'd283 && y == 203) || (x == 420 && y == 608) ||
		(x == 389 && y == 265) || (x == 7'd586 && y == 7'd551) || (x == 390 && y == 566) ||
		(x == 203 && y == 131) || (x == 7'd347 && y == 327) || (x == 7'd406 && y == 7'd429) ||
		(x == 7'd627 && y == 267) || (x == 7'd286 && y == 7'd271) || (x == 515 && y == 7'd431) ||
		(x == 7'd541 && y == 7'd399) || (x == 462 && y == 357) || (x == 7'd211 && y == 7'd122) ||
		(x == 7'd273 && y == 7'd280) || (x == 228 && y == 352) || (x == 7'd605 && y == 317) ||
		(x == 134 && y == 397) || (x == 7'd99 && y == 7'd563) || (x == 582 && y == 145) ||
		(x == 7'd301 && y == 7'd133) || (x == 431 && y == 541) || (x == 7'd190 && y == 7'd214) ||
		(x == 7'd427 && y == 7'd410) || (x == 314 && y == 608) || (x == 7'd237 && y == 5) ||
		(x == 7'd24 && y == 586) || (x == 7'd219 && y == 7'd309) || (x == 7'd441 && y == 7'd634) ||
		(x == 92 && y == 7'd11) || (x == 7'd515 && y == 7'd583) || (x == 7'd153 && y == 7'd268) ||
		(x == 7'd177 && y == 7'd391) || (x == 7'd597 && y == 324) || (x == 7'd407 && y == 436) ||
		(x == 7'd608 && y == 7'd292) || (x == 193 && y == 7'd100) || (x == 7'd446 && y == 481) ||
		(x == 7'd158 && y == 7'd388) || (x == 628 && y == 7'd77) || (x == 475 && y == 7'd149) ||
		(x == 555 && y == 199) || (x == 7'd493 && y == 7'd17) || (x == 453 && y == 7'd107) ||
		(x == 7'd216 && y == 7'd537) || (x == 7'd516 && y == 555) || (x == 7'd400 && y == 7'd442) ||
		(x == 7'd247 && y == 7'd233) || (x == 387 && y == 7'd337) || (x == 7'd562 && y == 7'd269) ||
		(x == 7'd566 && y == 301) || (x == 205 && y == 7'd90) || (x == 559 && y == 7'd339) ||
		(x == 7'd232 && y == 522) || (x == 7'd429 && y == 7'd522) || (x == 7'd462 && y == 277) ||
		(x == 307 && y == 7'd397) || (x == 7'd282 && y == 7'd388) || (x == 7'd639 && y == 7'd614) ||
		(x == 213 && y == 196) || (x == 7'd209 && y == 7'd155) || (x == 7'd144 && y == 7'd528) ||
		(x == 378 && y == 7'd38) || (x == 7'd511 && y == 7'd236) || (x == 7'd35 && y == 194) ||
		(x == 7'd624 && y == 7'd578) || (x == 629 && y == 385) || (x == 7'd381 && y == 7'd590) ||
		(x == 377 && y == 7'd167) || (x == 7'd181 && y == 7'd271) || (x == 7'd146 && y == 7'd313) ||
		(x == 364 && y == 434) || (x == 7'd461 && y == 7'd340) || (x == 217 && y == 172) ||
		(x == 227 && y == 7'd250) || (x == 409 && y == 7'd502) || (x == 7'd142 && y == 456) ||
		(x == 493 && y == 507) || (x == 7'd361 && y == 7'd636) || (x == 7'd476 && y == 398) ||
		(x == 7'd200 && y == 7'd586) || (x == 7'd426 && y == 7'd164) || (x == 7'd273 && y == 7'd12) ||
		(x == 7'd628 && y == 7'd353) || (x == 553 && y == 7'd193) || (x == 197 && y == 453) ||
		(x == 7'd136 && y == 7'd515) || (x == 7'd518 && y == 7'd233) || (x == 7'd497 && y == 457) ||
		(x == 7'd379 && y == 7'd461) || (x == 315 && y == 7'd484) || (x == 7'd181 && y == 7'd157) ||
		(x == 7'd296 && y == 546) || (x == 545 && y == 609) || (x == 538 && y == 7'd208) ||
		(x == 290 && y == 7'd45) || (x == 7'd359 && y == 353) || (x == 7'd577 && y == 7'd341) ||
		(x == 610 && y == 248) || (x == 601 && y == 252) || (x == 7'd154 && y == 326) ||
		(x == 7'd511 && y == 7'd104) || (x == 7'd133 && y == 217) || (x == 7'd13 && y == 7'd317) ||
		(x == 363 && y == 464) || (x == 512 && y == 447) || (x == 7'd225 && y == 578) ||
		(x == 7'd489 && y == 7'd502) || (x == 7'd166 && y == 349) || (x == 317 && y == 7'd441) ||
		(x == 7'd434 && y == 7'd389) || (x == 7'd155 && y == 539) || (x == 7'd494 && y == 7'd129) ||
		(x == 7'd549 && y == 618) || (x == 453 && y == 201) || (x == 578 && y == 7'd72) ||
		(x == 7'd36 && y == 380) || (x == 420 && y == 133) || (x == 7'd243 && y == 7'd633) ||
		(x == 7'd468 && y == 263) || (x == 252 && y == 7'd28) || (x == 7'd377 && y == 7'd491) ||
		(x == 7'd321 && y == 259) || (x == 7'd255 && y == 7'd98) || (x == 219 && y == 552) ||
		(x == 113 && y == 7'd526) || (x == 488 && y == 607) || (x == 579 && y == 7'd103) ||
		(x == 152 && y == 7'd35) || (x == 183 && y == 7'd217) || (x == 7'd100 && y == 355) ||
		(x == 7'd453 && y == 7'd34) || (x == 334 && y == 7'd45) || (x == 276 && y == 260) ||
		(x == 202 && y == 220) || (x == 7'd458 && y == 309) || (x == 7'd189 && y == 432) ||
		(x == 7'd424 && y == 7'd121) || (x == 7'd613 && y == 7'd131) || (x == 634 && y == 443) ||
		(x == 127 && y == 7'd355) || (x == 7'd240 && y == 7'd243) || (x == 357 && y == 7'd565) ||
		(x == 7'd587 && y == 493) || (x == 576 && y == 7'd13) || (x == 7'd263 && y == 621) ||
		(x == 7'd84 && y == 186) || (x == 7'd578 && y == 7'd562) || (x == 7'd608 && y == 7'd623) ||
		(x == 429 && y == 583) || (x == 558 && y == 607) || (x == 7'd538 && y == 621) ||
		(x == 633 && y == 7'd210) || (x == 311 && y == 7'd6) || (x == 504 && y == 7'd202) ||
		(x == 401 && y == 7'd257) || (x == 269 && y == 7'd442) || (x == 251 && y == 7'd310) ||
		(x == 88 && y == 81) || (x == 472 && y == 411) || (x == 7'd219 && y == 566) ||
		(x == 159 && y == 618) || (x == 7'd424 && y == 7'd340) || (x == 7'd452 && y == 7'd564) ||
		(x == 550 && y == 7'd287) || (x == 7'd127 && y == 179) || (x == 7'd542 && y == 600) ||
		(x == 7'd478 && y == 7'd397) || (x == 300 && y == 245) || (x == 7'd254 && y == 45) ||
		(x == 7'd515 && y == 317) || (x == 7'd16 && y == 7'd238) || (x == 178 && y == 7'd6) ||
		(x == 7'd376 && y == 627) || (x == 349 && y == 373) || (x == 500 && y == 267) ||
		(x == 7'd118 && y == 486) || (x == 7'd472 && y == 7'd551) || (x == 7'd186 && y == 170) ||
		(x == 7'd599 && y == 7'd373) || (x == 7'd405 && y == 395) || (x == 7'd231 && y == 262) ||
		(x == 7'd420 && y == 7'd448) || (x == 7'd598 && y == 558) || (x == 7'd425 && y == 7'd436) ||
		(x == 7'd274 && y == 510) || (x == 7'd264 && y == 7'd249) || (x == 7'd62 && y == 7'd340) ||
		(x == 7'd9 && y == 258) || (x == 584 && y == 7'd560) || (x == 7'd603 && y == 619) ||
		(x == 305 && y == 7'd218) || (x == 7'd457 && y == 271) || (x == 7'd102 && y == 580) ||
		(x == 400 && y == 372) || (x == 617 && y == 636) || (x == 458 && y == 288) ||
		(x == 7'd194 && y == 337) || (x == 7'd393 && y == 7'd279) || (x == 7'd538 && y == 7'd548) ||
		(x == 285 && y == 7'd240) || (x == 253 && y == 519) || (x == 232 && y == 7'd361) ||
		(x == 318 && y == 7'd43) || (x == 7'd320 && y == 116) || (x == 7'd251 && y == 7'd614) ||
		(x == 98 && y == 7'd169) || (x == 7'd302 && y == 176) || (x == 433 && y == 7'd270) ||
		(x == 7'd378 && y == 31) || (x == 380 && y == 7'd515) || (x == 7'd322 && y == 7'd219) ||
		(x == 7'd179 && y == 553) || (x == 7'd562 && y == 285) || (x == 563 && y == 520) ||
		(x == 7'd350 && y == 7'd163) || (x == 7'd313 && y == 7'd622) || (x == 7'd559 && y == 7'd516) ||
		(x == 7'd502 && y == 7'd549) || (x == 7'd530 && y == 7'd41) || (x == 433 && y == 7'd557) ||
		(x == 7'd160 && y == 239) || (x == 122 && y == 7'd261) || (x == 7'd484 && y == 501) ||
		(x == 443 && y == 7'd74) || (x == 7'd36 && y == 321) || (x == 7'd409 && y == 7'd636) ||
		(x == 7'd8 && y == 361) || (x == 606 && y == 239) || (x == 7'd314 && y == 7'd315) ||
		(x == 7'd14 && y == 587) || (x == 7'd206 && y == 223) || (x == 284 && y == 230) ||
		(x == 405 && y == 497) || (x == 7'd450 && y == 7'd502) || (x == 7'd240 && y == 7'd454) ||
		(x == 521 && y == 7'd105) || (x == 7'd552 && y == 143) || (x == 7'd362 && y == 7'd502) ||
		(x == 169 && y == 309) || (x == 4 && y == 7'd504) || (x == 7'd420 && y == 7'd403) ||
		(x == 7'd116 && y == 7'd380) || (x == 7'd624 && y == 632) || (x == 475 && y == 250) ||
		(x == 583 && y == 449) || (x == 7'd284 && y == 7'd432) || (x == 7'd265 && y == 7'd32) ||
		(x == 461 && y == 7'd126) || (x == 7'd478 && y == 7'd566) || (x == 207 && y == 159) ||
		(x == 410 && y == 147) || (x == 426 && y == 590) || (x == 7'd534 && y == 7'd415) ||
		(x == 7'd178 && y == 626) || (x == 7'd274 && y == 396) || (x == 7'd63 && y == 379) ||
		(x == 7'd386 && y == 7'd176) || (x == 340 && y == 7'd139) || (x == 2 && y == 7'd305) ||
		(x == 7'd431 && y == 296) || (x == 7'd441 && y == 7'd148) || (x == 7'd38 && y == 485) ||
		(x == 347 && y == 146) || (x == 397 && y == 7'd247) || (x == 7'd251 && y == 7'd567) ||
		(x == 193 && y == 7'd207) || (x == 7'd174 && y == 7'd264) || (x == 571 && y == 7'd639) ||
		(x == 488 && y == 631) || (x == 238 && y == 340) || (x == 7'd261 && y == 7'd610) ||
		(x == 7'd574 && y == 425) || (x == 497 && y == 7'd301) || (x == 7'd578 && y == 7'd61) ||
		(x == 345 && y == 541) || (x == 102 && y == 7'd462) || (x == 212 && y == 455) ||
		(x == 7'd379 && y == 7'd513) || (x == 7'd197 && y == 7'd461) || (x == 632 && y == 7'd159) ||
		(x == 7'd370 && y == 7'd67) || (x == 431 && y == 7'd128) || (x == 7'd450 && y == 7'd89) ||
		(x == 7'd168 && y == 553) || (x == 194 && y == 638) || (x == 7'd499 && y == 460) ||
		(x == 7'd373 && y == 624) || (x == 329 && y == 488) || (x == 7'd216 && y == 7'd147) ||
		(x == 441 && y == 7'd1) || (x == 495 && y == 507) || (x == 7'd7 && y == 7'd205) ||
		(x == 537 && y == 481) || (x == 7'd236 && y == 7'd244) || (x == 417 && y == 247) ||
		(x == 263 && y == 130) || (x == 302 && y == 356) || (x == 7'd113 && y == 7'd576) ||
		(x == 7'd289 && y == 304) || (x == 621 && y == 7'd243) || (x == 7'd473 && y == 120) ||
		(x == 7'd588 && y == 7'd415) || (x == 7'd567 && y == 138) || (x == 7'd289 && y == 635) ||
		(x == 636 && y == 7'd40) || (x == 7'd581 && y == 7'd181) || (x == 531 && y == 238) ||
		(x == 7'd468 && y == 609) || (x == 7'd331 && y == 310) || (x == 7'd204 && y == 248) ||
		(x == 7'd288 && y == 609) || (x == 7'd185 && y == 7'd595) || (x == 7'd346 && y == 7'd380) ||
		(x == 381 && y == 161) || (x == 18 && y == 7'd298) || (x == 7'd139 && y == 7'd164) ||
		(x == 7'd23 && y == 302) || (x == 535 && y == 7'd391) || (x == 400 && y == 7'd86) ||
		(x == 7'd319 && y == 583) || (x == 482 && y == 7'd629) || (x == 7'd457 && y == 616) ||
		(x == 205 && y == 7'd33) || (x == 151 && y == 7'd617) || (x == 7'd225 && y == 292) ||
		(x == 398 && y == 527) || (x == 7'd324 && y == 192) || (x == 17 && y == 7'd290) ||
		(x == 515 && y == 7'd130) || (x == 325 && y == 7'd43) || (x == 7'd350 && y == 7'd539) ||
		(x == 513 && y == 552) || (x == 7'd236 && y == 7'd503) || (x == 7'd441 && y == 7'd603) ||
		(x == 7'd493 && y == 51) || (x == 340 && y == 7'd245) || (x == 7'd446 && y == 7'd245) ||
		(x == 413 && y == 7'd577) || (x == 489 && y == 612) || (x == 149 && y == 7'd128) ||
		(x == 7'd91 && y == 7'd167) || (x == 370 && y == 7'd527) || (x == 7'd484 && y == 80) ||
		(x == 7'd238 && y == 7'd282) || (x == 7'd516 && y == 301) || (x == 7'd602 && y == 7'd228) ||
		(x == 7'd521 && y == 7'd244) || (x == 494 && y == 602) || (x == 7'd479 && y == 34) ||
		(x == 7'd6 && y == 7'd448) || (x == 7'd446 && y == 7'd138) || (x == 7'd112 && y == 7'd181) ||
		(x == 125 && y == 7'd249) || (x == 7'd445 && y == 7'd320) || (x == 271 && y == 7'd214) ||
		(x == 391 && y == 273) || (x == 7'd461 && y == 467) || (x == 178 && y == 541) ||
		(x == 7'd619 && y == 7'd506) || (x == 7'd459 && y == 7'd174) || (x == 23 && y == 7'd377) ||
		(x == 495 && y == 7'd208) || (x == 257 && y == 284) || (x == 7'd512 && y == 588) ||
		(x == 7'd516 && y == 7'd184) || (x == 515 && y == 7'd93) || (x == 7'd154 && y == 7'd156) ||
		(x == 7'd188 && y == 371) || (x == 7'd518 && y == 69) || (x == 7'd462 && y == 7'd220) ||
		(x == 504 && y == 571) || (x == 7'd605 && y == 181) || (x == 7'd290 && y == 88) ||
		(x == 7'd382 && y == 7'd144) || (x == 7'd314 && y == 14) || (x == 7'd506 && y == 61) ||
		(x == 278 && y == 7'd47) || (x == 7'd297 && y == 232) || (x == 7'd40 && y == 7'd378) ||
		(x == 552 && y == 7'd7) || (x == 7'd103 && y == 174) || (x == 7'd605 && y == 7'd520) ||
		(x == 279 && y == 7'd141) || (x == 7'd244 && y == 141) || (x == 462 && y == 7'd306) ||
		(x == 7'd312 && y == 7'd107) || (x == 411 && y == 477) || (x == 7'd17 && y == 7'd243) ||
		(x == 7'd9 && y == 7'd422) || (x == 7'd426 && y == 576) || (x == 451 && y == 278) ||
		(x == 7'd520 && y == 65) || (x == 482 && y == 7'd365) || (x == 233 && y == 7'd297) ||
		(x == 7'd302 && y == 539) || (x == 7'd606 && y == 508) || (x == 7'd406 && y == 7'd160) ||
		(x == 7'd574 && y == 7'd296) || (x == 7'd441 && y == 7'd71) || (x == 7'd262 && y == 7'd289) ||
		(x == 7'd67 && y == 7'd60) || (x == 7'd395 && y == 7'd80) || (x == 491 && y == 638) ||
		(x == 7'd350 && y == 7'd267) || (x == 7'd175 && y == 7'd202) || (x == 7'd533 && y == 79) ||
		(x == 7'd372 && y == 7'd546) || (x == 473 && y == 298) || (x == 147 && y == 455) ||
		(x == 262 && y == 389) || (x == 7'd498 && y == 53) || (x == 7'd524 && y == 479) ||
		(x == 7'd479 && y == 7'd366) || (x == 392 && y == 582) || (x == 7'd232 && y == 110) ||
		(x == 379 && y == 297) || (x == 121 && y == 7'd481) || (x == 551 && y == 132) ||
		(x == 332 && y == 7'd209) || (x == 188 && y == 7'd496) || (x == 634 && y == 7'd549) ||
		(x == 7'd391 && y == 516) || (x == 7'd137 && y == 7'd248) || (x == 7'd504 && y == 7'd425) ||
		(x == 402 && y == 415) || (x == 7'd638 && y == 438) || (x == 240 && y == 276) ||
		(x == 622 && y == 7'd559) || (x == 403 && y == 147) || (x == 7'd385 && y == 348) ||
		(x == 7'd552 && y == 7'd117) || (x == 7'd518 && y == 7'd249) || (x == 7'd267 && y == 224) ||
		(x == 7'd629 && y == 7'd329) || (x == 7'd505 && y == 371) || (x == 7'd503 && y == 266) ||
		(x == 7'd506 && y == 434) || (x == 313 && y == 596) || (x == 7'd227 && y == 7'd583) ||
		(x == 7'd100 && y == 355) || (x == 171 && y == 7'd541) || (x == 7'd475 && y == 7'd397) ||
		(x == 7'd11 && y == 366) || (x == 347 && y == 457) || (x == 7'd156 && y == 417) ||
		(x == 384 && y == 7'd484) || (x == 7'd456 && y == 582) || (x == 285 && y == 7'd47) ||
		(x == 412 && y == 7'd328) || (x == 7'd490 && y == 7'd148) || (x == 133 && y == 178) ||
		(x == 7'd321 && y == 7'd84) || (x == 5 && y == 7'd104) || (x == 562 && y == 7'd592) ||
		(x == 7'd331 && y == 259) || (x == 7'd498 && y == 7'd474) || (x == 100 && y == 7'd146) ||
		(x == 361 && y == 295) || (x == 511 && y == 348) || (x == 7'd540 && y == 390) ||
		(x == 272 && y == 7'd581) || (x == 217 && y == 390) || (x == 7'd122 && y == 7'd449) ||
		(x == 7'd422 && y == 7'd610) || (x == 7'd67 && y == 7'd390) || (x == 588 && y == 7'd138) ||
		(x == 7'd506 && y == 7'd142) || (x == 208 && y == 430) || (x == 7'd414 && y == 415) ||
		(x == 7'd529 && y == 473) || (x == 290 && y == 7'd132) || (x == 7'd230 && y == 7'd533) ||
		(x == 7'd354 && y == 7'd334) || (x == 442 && y == 7'd259) || (x == 186 && y == 480) ||
		(x == 531 && y == 317) || (x == 7'd55 && y == 471) || (x == 7'd630 && y == 7'd224) ||
		(x == 537 && y == 7'd208) || (x == 7'd254 && y == 7'd407) || (x == 7'd72 && y == 353) ||
		(x == 519 && y == 7'd459) || (x == 530 && y == 7'd498) || (x == 7'd233 && y == 375) ||
		(x == 7'd324 && y == 7'd595) || (x == 7'd298 && y == 7'd410) || (x == 7'd438 && y == 318) ||
		(x == 306 && y == 7'd8) || (x == 7'd474 && y == 7'd211) || (x == 195 && y == 7'd534) ||
		(x == 141 && y == 7'd297) || (x == 129 && y == 152) || (x == 7'd164 && y == 380) ||
		(x == 438 && y == 199) || (x == 202 && y == 7'd465) || (x == 7'd537 && y == 410) ||
		(x == 7'd550 && y == 198) || (x == 638 && y == 7'd551) || (x == 7'd161 && y == 7'd319) ||
		(x == 7'd198 && y == 371) || (x == 7'd403 && y == 65) || (x == 7'd363 && y == 7'd531) ||
		(x == 7'd363 && y == 7'd479) || (x == 535 && y == 594) || (x == 330 && y == 7'd100) ||
		(x == 489 && y == 192) || (x == 369 && y == 7'd536) || (x == 189 && y == 7'd151) ||
		(x == 7'd9 && y == 258) || (x == 461 && y == 7'd519) || (x == 373 && y == 589) ||
		(x == 7'd292 && y == 7'd443) || (x == 7'd401 && y == 83) || (x == 7'd61 && y == 244) ||
		(x == 7'd482 && y == 205) || (x == 7'd505 && y == 236) || (x == 7'd507 && y == 358) ||
		(x == 7'd160 && y == 171) || (x == 542 && y == 7'd6) || (x == 7'd437 && y == 201) ||
		(x == 256 && y == 566) || (x == 240 && y == 179) || (x == 7'd553 && y == 39) ||
		(x == 7'd435 && y == 461) || (x == 540 && y == 7'd121) || (x == 7'd78 && y == 613) ||
		(x == 130 && y == 7'd252) || (x == 23 && y == 122) || (x == 588 && y == 7'd3) ||
		(x == 467 && y == 7'd25) || (x == 7'd156 && y == 326) || (x == 7'd559 && y == 7'd541) ||
		(x == 348 && y == 382) || (x == 7'd260 && y == 154) || (x == 7'd640 && y == 317) ||
		(x == 7'd485 && y == 7'd391) || (x == 7'd552 && y == 7'd390) || (x == 615 && y == 331) ||
		(x == 496 && y == 7'd54) || (x == 7'd196 && y == 149) || (x == 7'd337 && y == 7'd637) ||
		(x == 408 && y == 7'd339) || (x == 275 && y == 7'd248) || (x == 326 && y == 264) ||
		(x == 7'd452 && y == 112) || (x == 71 && y == 7'd283) || (x == 618 && y == 7'd253) ||
		(x == 7'd263 && y == 453) || (x == 269 && y == 7'd126) || (x == 390 && y == 7'd422) ||
		(x == 7'd320 && y == 38) || (x == 7'd537 && y == 477) || (x == 7'd628 && y == 7'd92) ||
		(x == 7'd330 && y == 7'd1) || (x == 7'd565 && y == 572) || (x == 152 && y == 7'd152) ||
		(x == 7'd389 && y == 7'd10) || (x == 7'd362 && y == 7'd368) || (x == 7'd224 && y == 7'd492) ||
		(x == 148 && y == 7'd543) || (x == 7'd255 && y == 7'd242) || (x == 426 && y == 507) ||
		(x == 7'd250 && y == 287) || (x == 7'd500 && y == 7'd87) || (x == 239 && y == 512) ||
		(x == 7'd258 && y == 7'd10) || (x == 7'd569 && y == 166) || (x == 587 && y == 7'd223) ||
		(x == 623 && y == 7'd284) || (x == 7'd536 && y == 7'd431) || (x == 7'd404 && y == 69) ||
		(x == 171 && y == 7'd555) || (x == 392 && y == 235) || (x == 7'd255 && y == 7'd386) ||
		(x == 7'd506 && y == 7'd592) || (x == 7'd458 && y == 469) || (x == 7'd461 && y == 7'd179) ||
		(x == 398 && y == 238) || (x == 7'd139 && y == 7'd205) || (x == 487 && y == 187) ||
		(x == 185 && y == 280) || (x == 7'd125 && y == 163) || (x == 7'd454 && y == 489) ||
		(x == 7'd301 && y == 7'd357) || (x == 465 && y == 7'd534) || (x == 7'd500 && y == 151) ||
		(x == 592 && y == 221) || (x == 403 && y == 614) || (x == 7'd146 && y == 7'd578) ||
		(x == 224 && y == 7'd518) || (x == 268 && y == 406) || (x == 193 && y == 516) ||
		(x == 258 && y == 452) || (x == 372 && y == 361) || (x == 532 && y == 271) ||
		(x == 7'd595 && y == 7'd76) || (x == 596 && y == 7'd15) || (x == 238 && y == 468) ||
		(x == 7'd596 && y == 7'd414) || (x == 7'd469 && y == 605) || (x == 505 && y == 7'd398) ||
		(x == 519 && y == 530) || (x == 7'd579 && y == 7'd211) || (x == 254 && y == 7'd463) ||
		(x == 7'd410 && y == 426) || (x == 7'd325 && y == 7'd572) || (x == 320 && y == 571) ||
		(x == 566 && y == 434) || (x == 7'd178 && y == 613) || (x == 573 && y == 7'd362) ||
		(x == 7'd454 && y == 7'd561) || (x == 7'd315 && y == 7'd247) || (x == 7'd70 && y == 7'd522) ||
		(x == 7'd165 && y == 7'd598) || (x == 7'd135 && y == 7'd458) || (x == 345 && y == 7'd573) ||
		(x == 7'd346 && y == 7'd164) || (x == 77 && y == 7'd542) || (x == 340 && y == 134) ||
		(x == 191 && y == 185) || (x == 7'd46 && y == 7'd526) || (x == 406 && y == 7'd71) ||
		(x == 443 && y == 450) || (x == 7'd563 && y == 404) || (x == 193 && y == 465) ||
		(x == 278 && y == 540) || (x == 127 && y == 7'd458) || (x == 7'd126 && y == 7'd297) ||
		(x == 7'd165 && y == 7'd241) || (x == 183 && y == 332) || (x == 7'd548 && y == 107) ||
		(x == 300 && y == 443) || (x == 391 && y == 465) || (x == 7'd254 && y == 534) ||
		(x == 7'd134 && y == 7'd223) || (x == 7'd115 && y == 7'd194) || (x == 404 && y == 7'd54) ||
		(x == 379 && y == 7'd71) || (x == 7'd109 && y == 565) || (x == 7'd490 && y == 522) ||
		(x == 7'd106 && y == 100) || (x == 169 && y == 130) || (x == 572 && y == 7'd539) ||
		(x == 311 && y == 7'd480) || (x == 7'd468 && y == 445) || (x == 7'd317 && y == 7'd473) ||
		(x == 7'd494 && y == 7'd168) || (x == 629 && y == 333) || (x == 7'd484 && y == 7'd178) ||
		(x == 346 && y == 242) || (x == 234 && y == 333) || (x == 7'd324 && y == 571) ||
		(x == 7'd77 && y == 7'd380) || (x == 7'd309 && y == 512) || (x == 7'd287 && y == 358) ||
		(x == 7'd629 && y == 7'd381) || (x == 7'd211 && y == 7'd447) || (x == 7'd484 && y == 7'd229) ||
		(x == 246 && y == 7'd286) || (x == 7'd474 && y == 7'd522) || (x == 286 && y == 357) ||
		(x == 7'd276 && y == 7'd270) || (x == 118 && y == 7'd415) || (x == 7'd344 && y == 134) ||
		(x == 524 && y == 529) || (x == 256 && y == 7'd236) || (x == 218 && y == 165) ||
		(x == 7'd249 && y == 7'd289) || (x == 7'd470 && y == 7'd436) || (x == 7'd454 && y == 220) ||
		(x == 244 && y == 7'd521) || (x == 7'd545 && y == 7'd144) || (x == 494 && y == 7'd359) ||
		(x == 516 && y == 254) || (x == 7'd268 && y == 22) || (x == 7'd503 && y == 7'd423) ||
		(x == 7'd304 && y == 230) || (x == 7'd280 && y == 380) || (x == 14 && y == 7'd569) ||
		(x == 93 && y == 7'd463) || (x == 7'd21 && y == 376) || (x == 7'd433 && y == 581) ||
		(x == 7'd628 && y == 7'd141) || (x == 420 && y == 201) || (x == 7'd211 && y == 7'd65) ||
		(x == 578 && y == 162) || (x == 569 && y == 7'd328) || (x == 516 && y == 7'd168) ||
		(x == 21 && y == 7'd582) || (x == 7'd69 && y == 7'd294) || (x == 7'd154 && y == 7'd558) ||
		(x == 7'd396 && y == 296) || (x == 7'd122 && y == 7'd248) || (x == 7'd595 && y == 290) ||
		(x == 497 && y == 403) || (x == 7'd289 && y == 7'd313) || (x == 7'd267 && y == 44) ||
		(x == 616 && y == 7'd279) || (x == 7'd543 && y == 7'd587) || (x == 7'd286 && y == 7'd579) ||
		(x == 7'd639 && y == 135) || (x == 7'd625 && y == 596) || (x == 7'd346 && y == 433) ||
		(x == 391 && y == 7'd181) || (x == 7'd495 && y == 7'd528) || (x == 169 && y == 7'd251) ||
		(x == 91 && y == 7'd496) || (x == 7'd310 && y == 7'd406) || (x == 7'd267 && y == 433) ||
		(x == 7'd573 && y == 7'd628) || (x == 7'd522 && y == 278) || (x == 545 && y == 7'd196) ||
		(x == 7'd337 && y == 7'd153) || (x == 372 && y == 7'd84) || (x == 588 && y == 7'd482) ||
		(x == 7'd45 && y == 598) || (x == 163 && y == 7'd383) || (x == 40 && y == 7'd15) ||
		(x == 7'd404 && y == 7'd635) || (x == 7'd211 && y == 7'd208) || (x == 99 && y == 7'd492) ||
		(x == 7'd569 && y == 267) || (x == 487 && y == 7'd515) || (x == 490 && y == 535) ||
		(x == 7'd499 && y == 535) || (x == 408 && y == 7'd80) || (x == 422 && y == 550) ||
		(x == 400 && y == 7'd502) || (x == 360 && y == 244) || (x == 210 && y == 7'd85) ||
		(x == 7'd71 && y == 124) || (x == 476 && y == 7'd460) || (x == 7'd109 && y == 7'd560) ||
		(x == 7'd192 && y == 466) || (x == 194 && y == 353) || (x == 7'd603 && y == 7'd625) ||
		(x == 7'd66 && y == 57) || (x == 7'd423 && y == 518) || (x == 472 && y == 292) ||
		(x == 7'd474 && y == 199) || (x == 7'd635 && y == 7'd380) || (x == 189 && y == 294) ||
		(x == 7'd189 && y == 7'd301) || (x == 391 && y == 484) || (x == 7'd104 && y == 522) ||
		(x == 466 && y == 7'd250) || (x == 7'd35 && y == 499) || (x == 7'd172 && y == 303) ||
		(x == 7'd404 && y == 603) || (x == 507 && y == 382) || (x == 7'd50 && y == 439) ||
		(x == 129 && y == 598) || (x == 7'd184 && y == 521) || (x == 7'd104 && y == 7'd431) ||
		(x == 7'd493 && y == 7'd114) || (x == 7'd520 && y == 7'd149) || (x == 633 && y == 7'd406) ||
		(x == 520 && y == 7'd139) || (x == 374 && y == 633) || (x == 605 && y == 7'd85) ||
		(x == 7'd257 && y == 244) || (x == 590 && y == 7'd123) || (x == 7'd377 && y == 7'd485) ||
		(x == 7'd196 && y == 7'd100) || (x == 349 && y == 480) || (x == 7'd135 && y == 7'd453) ||
		(x == 7'd361 && y == 355) || (x == 534 && y == 284) || (x == 190 && y == 228) ||
		(x == 7'd445 && y == 7'd523) || (x == 7'd357 && y == 401) || (x == 7'd74 && y == 372) ||
		(x == 139 && y == 7'd573) || (x == 132 && y == 7'd632) || (x == 7'd157 && y == 7'd385) ||
		(x == 7'd127 && y == 308) || (x == 632 && y == 481) || (x == 156 && y == 639) ||
		(x == 330 && y == 405) || (x == 7'd630 && y == 7'd266) || (x == 219 && y == 461) ||
		(x == 182 && y == 7'd192) || (x == 7'd180 && y == 7'd130) || (x == 7'd379 && y == 144) ||
		(x == 342 && y == 7'd247) || (x == 360 && y == 220) || (x == 7'd608 && y == 7'd468) ||
		(x == 7'd545 && y == 7'd466) || (x == 576 && y == 580) || (x == 377 && y == 7'd368) ||
		(x == 270 && y == 452) || (x == 66 && y == 7'd187) || (x == 7'd293 && y == 7'd341) ||
		(x == 7'd624 && y == 634) || (x == 298 && y == 496) || (x == 7'd526 && y == 7'd598) ||
		(x == 147 && y == 358) || (x == 7'd197 && y == 630) || (x == 475 && y == 7'd51) ||
		(x == 633 && y == 7'd602) || (x == 516 && y == 573) || (x == 589 && y == 7'd638) ||
		(x == 416 && y == 413) || (x == 7'd212 && y == 7'd333) || (x == 7'd608 && y == 7'd435) ||
		(x == 390 && y == 496) || (x == 7'd439 && y == 7'd324) || (x == 431 && y == 7'd256) ||
		(x == 160 && y == 7'd111) || (x == 195 && y == 531) || (x == 7'd64 && y == 457) ||
		(x == 439 && y == 7'd608) || (x == 7'd363 && y == 220) || (x == 379 && y == 7'd359) ||
		(x == 7'd448 && y == 7'd88) || (x == 7'd481 && y == 413) || (x == 213 && y == 235) ||
		(x == 7'd308 && y == 302) || (x == 243 && y == 7'd441) || (x == 7'd21 && y == 530) ||
		(x == 7'd8 && y == 524) || (x == 7'd488 && y == 7'd484) || (x == 7'd621 && y == 7'd412) ||
		(x == 7'd221 && y == 7'd164) || (x == 7'd351 && y == 471) || (x == 7'd494 && y == 7'd413) ||
		(x == 7'd613 && y == 7'd336) || (x == 7'd249 && y == 7'd518) || (x == 7'd18 && y == 333) ||
		(x == 562 && y == 314) || (x == 180 && y == 502) || (x == 147 && y == 7'd515) ||
		(x == 7'd38 && y == 7'd129) || (x == 504 && y == 600) || (x == 262 && y == 7'd370) ||
		(x == 7'd625 && y == 248) || (x == 7'd404 && y == 7'd506) || (x == 7'd615 && y == 7'd297) ||
		(x == 306 && y == 7'd394) || (x == 339 && y == 7'd437) || (x == 7'd10 && y == 7'd162) ||
		(x == 7'd485 && y == 7'd105) || (x == 7'd612 && y == 296) || (x == 7'd534 && y == 372) ||
		(x == 7'd522 && y == 78) || (x == 7'd630 && y == 7'd314) || (x == 7'd323 && y == 259) ||
		(x == 7'd67 && y == 7'd635) || (x == 7'd313 && y == 514) || (x == 168 && y == 135) ||
		(x == 7'd392 && y == 15) || (x == 283 && y == 465) || (x == 224 && y == 570) ||
		(x == 178 && y == 7'd261) || (x == 433 && y == 246) || (x == 7'd269 && y == 7'd496) ||
		(x == 7'd80 && y == 253) || (x == 7'd267 && y == 7'd404) || (x == 7'd403 && y == 7'd266) ||
		(x == 7'd503 && y == 7'd389) || (x == 518 && y == 7'd549) || (x == 7'd474 && y == 204) ||
		(x == 335 && y == 7'd491) || (x == 468 && y == 7'd1) || (x == 531 && y == 7'd63) ||
		(x == 7'd464 && y == 490) || (x == 7'd609 && y == 7'd237) || (x == 312 && y == 468) ||
		(x == 131 && y == 7'd535) || (x == 7'd467 && y == 7'd327) || (x == 7'd511 && y == 430) ||
		(x == 7'd243 && y == 589) || (x == 7'd139 && y == 111) || (x == 342 && y == 7'd297) ||
		(x == 7'd520 && y == 7'd77) || (x == 219 && y == 7'd186) || (x == 149 && y == 7'd606) ||
		(x == 406 && y == 600) || (x == 7'd104 && y == 217) || (x == 552 && y == 480) ||
		(x == 7'd48 && y == 7'd361) || (x == 221 && y == 621) || (x == 366 && y == 548) ||
		(x == 7'd387 && y == 7'd198) || (x == 7'd223 && y == 7'd392) || (x == 7'd285 && y == 337) ||
		(x == 7'd381 && y == 183) || (x == 7'd629 && y == 7'd597) || (x == 7'd473 && y == 294) ||
		(x == 7'd392 && y == 366) || (x == 7'd407 && y == 7'd559) || (x == 410 && y == 535) ||
		(x == 590 && y == 209) || (x == 7'd496 && y == 7'd268) || (x == 257 && y == 7'd430) ||
		(x == 608 && y == 223) || (x == 251 && y == 577) || (x == 577 && y == 7'd196) ||
		(x == 7'd454 && y == 499) || (x == 265 && y == 289) || (x == 7'd573 && y == 7'd579) ||
		(x == 7'd633 && y == 7'd376) || (x == 7'd63 && y == 283) || (x == 7'd632 && y == 7'd85) ||
		(x == 405 && y == 7'd582) || (x == 388 && y == 562) || (x == 359 && y == 508) ||
		(x == 7'd471 && y == 305) || (x == 7'd144 && y == 414) || (x == 571 && y == 7'd417) ||
		(x == 41 && y == 7'd522) || (x == 323 && y == 251) || (x == 7'd12 && y == 7'd529) ||
		(x == 332 && y == 7'd379) || (x == 297 && y == 7'd389) || (x == 7'd394 && y == 7'd204) ||
		(x == 7'd11 && y == 154) || (x == 275 && y == 7'd252) || (x == 610 && y == 491) ||
		(x == 639 && y == 424) || (x == 7'd553 && y == 7'd263) || (x == 7'd83 && y == 7'd205) ||
		(x == 514 && y == 7'd111) || (x == 7'd509 && y == 7'd257) || (x == 29 && y == 7'd524) ||
		(x == 201 && y == 334) || (x == 7'd639 && y == 46) || (x == 166 && y == 464) ||
		(x == 7'd376 && y == 7'd548) || (x == 7'd299 && y == 530) || (x == 7'd480 && y == 412) ||
		(x == 7'd238 && y == 425) || (x == 7'd601 && y == 275) || (x == 144 && y == 271) ||
		(x == 290 && y == 505) || (x == 7'd362 && y == 120) || (x == 7'd158 && y == 2) ||
		(x == 222 && y == 7'd252) || (x == 7'd520 && y == 7'd500) || (x == 7'd324 && y == 637) ||
		(x == 7'd438 && y == 7'd494) || (x == 7'd635 && y == 7'd167) || (x == 7'd402 && y == 502) ||
		(x == 254 && y == 497) || (x == 7'd592 && y == 460) || (x == 412 && y == 369) ||
		(x == 7'd239 && y == 603) || (x == 7'd29 && y == 7'd302) || (x == 7'd258 && y == 7'd310) ||
		(x == 7'd37 && y == 7'd352) || (x == 191 && y == 7'd554) || (x == 7'd422 && y == 7'd584) ||
		(x == 170 && y == 7'd202) || (x == 546 && y == 416) || (x == 252 && y == 7'd207) ||
		(x == 7'd137 && y == 7'd426) || (x == 434 && y == 7'd66) || (x == 215 && y == 7'd175) ||
		(x == 7'd120 && y == 7'd621) || (x == 7'd155 && y == 7'd7) || (x == 7'd132 && y == 7'd200) ||
		(x == 7'd323 && y == 7'd636) || (x == 7'd443 && y == 7'd578) || (x == 7'd244 && y == 59) ||
		(x == 339 && y == 353) || (x == 7'd251 && y == 7'd189) || (x == 503 && y == 520) ||
		(x == 7'd421 && y == 205) || (x == 7'd3 && y == 336) || (x == 7'd545 && y == 7'd376) ||
		(x == 7'd14 && y == 246) || (x == 7'd577 && y == 7'd484) || (x == 7'd521 && y == 7'd368) ||
		(x == 7'd286 && y == 7'd481) || (x == 418 && y == 524) || (x == 7'd462 && y == 331) ||
		(x == 7'd196 && y == 7'd116) || (x == 7'd85 && y == 530) || (x == 418 && y == 7'd261) ||
		(x == 361 && y == 634) || (x == 364 && y == 381) || (x == 537 && y == 338) ||
		(x == 559 && y == 7'd625) || (x == 7'd580 && y == 7'd120) || (x == 312 && y == 7'd264) ||
		(x == 7'd348 && y == 7'd137) || (x == 473 && y == 7'd399) || (x == 7'd377 && y == 61) ||
		(x == 184 && y == 7'd241) || (x == 263 && y == 339) || (x == 7'd582 && y == 7'd179) ||
		(x == 7'd517 && y == 425) || (x == 7'd261 && y == 7'd290) || (x == 7'd430 && y == 7'd634) ||
		(x == 7'd588 && y == 7'd275) || (x == 7'd116 && y == 292) || (x == 7'd15 && y == 7'd400) ||
		(x == 366 && y == 491) || (x == 558 && y == 7'd365) || (x == 161 && y == 7'd392) ||
		(x == 130 && y == 7'd189) || (x == 7'd160 && y == 243) || (x == 7'd404 && y == 382) ||
		(x == 341 && y == 516) || (x == 634 && y == 487) || (x == 7'd605 && y == 7'd414) ||
		(x == 193 && y == 447) || (x == 436 && y == 555) || (x == 7'd216 && y == 7'd44) ||
		(x == 79 && y == 7'd595) || (x == 404 && y == 7'd145) || (x == 7'd635 && y == 53) ||
		(x == 7'd554 && y == 7'd8) || (x == 602 && y == 614) || (x == 7'd90 && y == 7'd181) ||
		(x == 351 && y == 7'd617) || (x == 7'd222 && y == 521) || (x == 7'd377 && y == 7'd519) ||
		(x == 7'd399 && y == 7'd60) || (x == 7'd201 && y == 7'd353) || (x == 7'd480 && y == 7'd266) ||
		(x == 7'd52 && y == 378) || (x == 338 && y == 253) || (x == 7'd15 && y == 142) ||
		(x == 7'd615 && y == 7'd276) || (x == 7'd441 && y == 7'd240) || (x == 7'd614 && y == 7'd311) ||
		(x == 7'd101 && y == 7'd488) || (x == 335 && y == 550) || (x == 7'd402 && y == 7'd321) ||
		(x == 7'd273 && y == 553) || (x == 262 && y == 376) || (x == 564 && y == 408) ||
		(x == 364 && y == 7'd403) || (x == 7'd111 && y == 358) || (x == 7'd351 && y == 9) ||
		(x == 7'd467 && y == 618) || (x == 7'd370 && y == 30) || (x == 7'd254 && y == 7'd540) ||
		(x == 7'd102 && y == 7'd557) || (x == 35 && y == 7'd498) || (x == 425 && y == 7'd404) ||
		(x == 491 && y == 7'd247) || (x == 7'd577 && y == 7'd582) || (x == 315 && y == 165) ||
		(x == 7'd487 && y == 7'd409) || (x == 7'd25 && y == 7'd434) || (x == 7'd636 && y == 7'd612) ||
		(x == 89 && y == 7'd175) || (x == 7'd475 && y == 7'd418) || (x == 7'd471 && y == 7'd300) ||
		(x == 7'd270 && y == 282) || (x == 429 && y == 7'd234) || (x == 7'd170 && y == 7'd153) ||
		(x == 204 && y == 203) || (x == 7'd143 && y == 115) || (x == 638 && y == 136) ||
		(x == 7'd396 && y == 7'd271) || (x == 143 && y == 341) || (x == 528 && y == 213) ||
		(x == 7'd539 && y == 145) || (x == 7'd276 && y == 7'd156) || (x == 7'd392 && y == 94) ||
		(x == 7'd16 && y == 310) || (x == 485 && y == 7'd455) || (x == 7'd608 && y == 565) ||
		(x == 621 && y == 7'd202) || (x == 550 && y == 7'd574) || (x == 138 && y == 7'd609) ||
		(x == 7'd523 && y == 18) || (x == 416 && y == 7'd394) || (x == 7'd66 && y == 637) ||
		(x == 7'd501 && y == 7'd107) || (x == 7'd325 && y == 329) || (x == 7'd567 && y == 7'd363) ||
		(x == 566 && y == 7'd73) || (x == 7'd559 && y == 7'd540) || (x == 7'd496 && y == 361) ||
		(x == 7'd395 && y == 412) || (x == 7'd242 && y == 7'd475) || (x == 611 && y == 299) ||
		(x == 7'd548 && y == 137) || (x == 154 && y == 7'd564) || (x == 7'd489 && y == 7'd111) ||
		(x == 633 && y == 563) || (x == 284 && y == 372) || (x == 7'd496 && y == 7'd242) ||
		(x == 89 && y == 7'd211) || (x == 7'd555 && y == 486) || (x == 392 && y == 395) ||
		(x == 393 && y == 7'd49) || (x == 7'd370 && y == 7'd287) || (x == 7'd251 && y == 7'd172) ||
		(x == 584 && y == 7'd576) || (x == 7'd418 && y == 7'd233) || (x == 7'd231 && y == 333) ||
		(x == 7'd207 && y == 7'd224) || (x == 7'd343 && y == 7'd207) || (x == 476 && y == 7'd391) ||
		(x == 7'd317 && y == 7'd283) || (x == 283 && y == 7'd135) || (x == 264 && y == 292) ||
		(x == 7'd392 && y == 7'd272) || (x == 7'd506 && y == 79) || (x == 7'd503 && y == 543) ||
		(x == 7'd340 && y == 7'd464) || (x == 458 && y == 520) || (x == 7'd368 && y == 7'd41) ||
		(x == 7'd378 && y == 7'd101) || (x == 7'd324 && y == 7'd233) || (x == 262 && y == 588) ||
		(x == 126 && y == 7'd81) || (x == 7'd91 && y == 452) || (x == 174 && y == 331) ||
		(x == 7'd211 && y == 406) || (x == 7'd588 && y == 7'd18) || (x == 577 && y == 244) ||
		(x == 7'd285 && y == 179) || (x == 297 && y == 7'd218) || (x == 346 && y == 7'd182) ||
		(x == 7'd472 && y == 637) || (x == 7'd165 && y == 7'd528) || (x == 7'd298 && y == 376) ||
		(x == 399 && y == 465) || (x == 7'd84 && y == 508) || (x == 7'd49 && y == 419) ||
		(x == 7'd276 && y == 7'd414) || (x == 7'd609 && y == 106) || (x == 7'd515 && y == 500) ||
		(x == 7'd116 && y == 155) || (x == 597 && y == 547) || (x == 122 && y == 7'd527) ||
		(x == 7'd529 && y == 7'd209) || (x == 7'd18 && y == 7'd195) || (x == 7'd477 && y == 7'd161) ||
		(x == 438 && y == 7'd553) || (x == 234 && y == 7'd373) || (x == 7'd206 && y == 7'd125) ||
		(x == 7'd217 && y == 449) || (x == 7'd487 && y == 7'd466) || (x == 630 && y == 7'd320) ||
		(x == 7'd579 && y == 7'd136) || (x == 7'd360 && y == 7'd633) || (x == 465 && y == 281) ||
		(x == 585 && y == 385) || (x == 7'd480 && y == 343) || (x == 7'd622 && y == 168) ||
		(x == 7'd44 && y == 184) || (x == 459 && y == 178) || (x == 7'd230 && y == 7'd562) ||
		(x == 490 && y == 7'd365) || (x == 258 && y == 7'd248) || (x == 7'd105 && y == 416) ||
		(x == 7'd594 && y == 7'd438) || (x == 7'd476 && y == 7'd160) || (x == 542 && y == 7'd229) ||
		(x == 443 && y == 197) || (x == 7'd140 && y == 553) || (x == 534 && y == 218) ||
		(x == 7'd524 && y == 263) || (x == 238 && y == 7'd586) || (x == 451 && y == 7'd322) ||
		(x == 7'd127 && y == 589) || (x == 504 && y == 343) || (x == 7'd523 && y == 7'd576) ||
		(x == 156 && y == 7'd147) || (x == 7'd464 && y == 140) || (x == 7'd373 && y == 7'd188) ||
		(x == 7'd204 && y == 7'd47) || (x == 133 && y == 305) || (x == 7'd399 && y == 7'd441) ||
		(x == 7'd573 && y == 377) || (x == 7'd282 && y == 254) || (x == 531 && y == 413) ||
		(x == 7'd68 && y == 7'd518) || (x == 432 && y == 264) || (x == 558 && y == 7'd366) ||
		(x == 160 && y == 7'd254) || (x == 421 && y == 286) || (x == 7'd474 && y == 469) ||
		(x == 7'd381 && y == 244) || (x == 358 && y == 7'd500) || (x == 364 && y == 7'd214) ||
		(x == 7'd532 && y == 7'd312) || (x == 322 && y == 7'd361) || (x == 473 && y == 7'd500) ||
		(x == 548 && y == 457) || (x == 7'd363 && y == 391) || (x == 7'd573 && y == 7'd471) ||
		(x == 197 && y == 7'd462) || (x == 31 && y == 7'd16) || (x == 7'd506 && y == 573) ||
		(x == 463 && y == 7'd281) || (x == 173 && y == 7'd585) || (x == 7'd375 && y == 62) ||
		(x == 7'd324 && y == 7'd524) || (x == 351 && y == 519) || (x == 7'd596 && y == 7'd257) ||
		(x == 439 && y == 7'd165) || (x == 7'd136 && y == 7'd630) || (x == 7'd531 && y == 7'd270) ||
		(x == 7'd434 && y == 7'd78) || (x == 266 && y == 254) || (x == 7'd129 && y == 429) ||
		(x == 7'd489 && y == 434) || (x == 279 && y == 593) || (x == 7'd176 && y == 7'd486) ||
		(x == 551 && y == 7'd224) || (x == 7'd296 && y == 7'd116) || (x == 639 && y == 592) ||
		(x == 229 && y == 150) || (x == 485 && y == 7'd333) || (x == 7'd136 && y == 7'd202) ||
		(x == 7'd412 && y == 7'd395) || (x == 7'd430 && y == 365) || (x == 7'd519 && y == 7'd310) ||
		(x == 109 && y == 7'd371) || (x == 445 && y == 7'd256) || (x == 7'd70 && y == 437) ||
		(x == 7'd96 && y == 340) || (x == 7'd107 && y == 7'd145) || (x == 201 && y == 7'd639) ||
		(x == 7'd30 && y == 7'd13) || (x == 7'd319 && y == 403) || (x == 7'd339 && y == 145) ||
		(x == 263 && y == 7'd407) || (x == 7'd332 && y == 7'd94) || (x == 278 && y == 525) ||
		(x == 7'd258 && y == 7'd411) || (x == 191 && y == 379) || (x == 7'd328 && y == 7'd253) ||
		(x == 7'd282 && y == 7'd459) || (x == 194 && y == 323) || (x == 7'd428 && y == 553) ||
		(x == 260 && y == 7'd351) || (x == 7'd574 && y == 581) || (x == 7'd189 && y == 7'd43) ||
		(x == 564 && y == 428) || (x == 7'd247 && y == 7'd340) || (x == 7'd220 && y == 423) ||
		(x == 446 && y == 7'd117) || (x == 174 && y == 228) || (x == 509 && y == 7'd94) ||
		(x == 223 && y == 609) || (x == 221 && y == 258) || (x == 247 && y == 7'd539) ||
		(x == 7'd405 && y == 7'd332) || (x == 7'd333 && y == 367) || (x == 7'd617 && y == 363) ||
		(x == 7'd134 && y == 468) || (x == 614 && y == 535) || (x == 280 && y == 7'd379) ||
		(x == 7'd360 && y == 569) || (x == 7'd373 && y == 7'd442) || (x == 120 && y == 7'd446) ||
		(x == 7'd367 && y == 7'd273) || (x == 7'd158 && y == 7'd385) || (x == 7'd608 && y == 261) ||
		(x == 7'd383 && y == 86) || (x == 192 && y == 307) || (x == 191 && y == 509) ||
		(x == 240 && y == 218) || (x == 7'd25 && y == 7'd510) || (x == 524 && y == 208) ||
		(x == 7'd543 && y == 7'd209) || (x == 7'd335 && y == 7'd432) || (x == 546 && y == 7'd170) ||
		(x == 7'd433 && y == 280) || (x == 209 && y == 275) || (x == 7'd137 && y == 7'd337) ||
		(x == 7'd331 && y == 7'd173) || (x == 283 && y == 7'd592) || (x == 92 && y == 7'd626) ||
		(x == 7'd633 && y == 457) || (x == 7'd444 && y == 7'd363) || (x == 190 && y == 375) ||
		(x == 393 && y == 7'd471) || (x == 92 && y == 7'd37) || (x == 457 && y == 7'd565) ||
		(x == 334 && y == 7'd399) || (x == 558 && y == 7'd178) || (x == 633 && y == 7'd347) ||
		(x == 7'd530 && y == 7'd516) || (x == 308 && y == 7'd197) || (x == 505 && y == 7'd332) ||
		(x == 271 && y == 7'd427) || (x == 7'd585 && y == 7'd554) || (x == 7'd29 && y == 7'd336) ||
		(x == 7'd570 && y == 7'd627) || (x == 95 && y == 7'd624) || (x == 132 && y == 626) ||
		(x == 7'd147 && y == 7'd582) || (x == 600 && y == 143) || (x == 7'd606 && y == 574) ||
		(x == 251 && y == 441) || (x == 7'd583 && y == 7'd298) || (x == 7'd111 && y == 243) ||
		(x == 7'd531 && y == 7'd327) || (x == 7'd593 && y == 319) || (x == 7'd424 && y == 479) ||
		(x == 293 && y == 451) || (x == 260 && y == 517) || (x == 540 && y == 134) ||
		(x == 100 && y == 7'd334) || (x == 171 && y == 7'd357) || (x == 3 && y == 7'd562) ||
		(x == 313 && y == 133) || (x == 476 && y == 7'd345) || (x == 7'd300 && y == 7'd134) ||
		(x == 7'd621 && y == 7'd153) || (x == 7'd347 && y == 114) || (x == 148 && y == 549) ||
		(x == 7'd320 && y == 637) || (x == 7'd337 && y == 7'd494) || (x == 326 && y == 619) ||
		(x == 7'd594 && y == 7'd564) || (x == 7'd573 && y == 33) || (x == 259 && y == 418) ||
		(x == 7'd32 && y == 7'd507) || (x == 7'd277 && y == 7'd287) || (x == 382 && y == 7'd495) ||
		(x == 8 && y == 45) || (x == 7'd231 && y == 232) || (x == 7'd122 && y == 7'd272) ||
		(x == 7'd262 && y == 7'd589) || (x == 548 && y == 421) || (x == 7'd168 && y == 7'd489) ||
		(x == 7'd550 && y == 7'd258) || (x == 7'd225 && y == 436) || (x == 7'd522 && y == 293) ||
		(x == 26 && y == 7'd268) || (x == 265 && y == 7'd164) || (x == 7'd290 && y == 7'd144) ||
		(x == 7'd9 && y == 179) || (x == 7'd598 && y == 607) || (x == 340 && y == 307) ||
		(x == 7'd539 && y == 7'd302) || (x == 7'd346 && y == 7'd355) || (x == 516 && y == 7'd594) ||
		(x == 7'd210 && y == 7'd178) || (x == 7'd403 && y == 561) || (x == 7'd429 && y == 7'd7) ||
		(x == 506 && y == 7'd390) || (x == 7'd348 && y == 141) || (x == 531 && y == 7'd292) ||
		(x == 7'd437 && y == 7'd279) || (x == 7'd155 && y == 7'd305) || (x == 7'd370 && y == 7'd635) ||
		(x == 211 && y == 7'd527) || (x == 7'd159 && y == 7'd387) || (x == 415 && y == 7'd26) ||
		(x == 7'd622 && y == 528) || (x == 174 && y == 540) || (x == 7'd268 && y == 7'd424) ||
		(x == 353 && y == 7'd455) || (x == 7'd268 && y == 19) || (x == 7'd239 && y == 7'd435) ||
		(x == 7'd411 && y == 7'd289) || (x == 7'd516 && y == 7'd27) || (x == 57 && y == 7'd86) ||
		(x == 463 && y == 511) || (x == 185 && y == 7'd213) || (x == 251 && y == 227) ||
		(x == 436 && y == 246) || (x == 313 && y == 7'd17) || (x == 7'd115 && y == 179) ||
		(x == 7'd383 && y == 7'd512) || (x == 7'd353 && y == 510) || (x == 295 && y == 7'd312) ||
		(x == 7'd234 && y == 7'd215) || (x == 169 && y == 7'd372) || (x == 345 && y == 7'd530) ||
		(x == 611 && y == 412) || (x == 556 && y == 7'd310) || (x == 7'd526 && y == 7'd56) ||
		(x == 7'd205 && y == 7'd148) || (x == 7'd282 && y == 7'd202) || (x == 248 && y == 251) ||
		(x == 7'd534 && y == 337) || (x == 7'd344 && y == 7'd166) || (x == 124 && y == 7'd335) ||
		(x == 7'd520 && y == 7'd62) || (x == 7'd559 && y == 435) || (x == 7'd69 && y == 576) ||
		(x == 538 && y == 512) || (x == 7'd506 && y == 7'd631) || (x == 7'd319 && y == 69) ||
		(x == 7'd395 && y == 34) || (x == 7'd263 && y == 31) || (x == 7'd632 && y == 7'd102) ||
		(x == 7'd216 && y == 624) || (x == 91 && y == 7'd89) || (x == 410 && y == 7'd472) ||
		(x == 511 && y == 345) || (x == 7'd241 && y == 570) || (x == 252 && y == 7'd299) ||
		(x == 7'd134 && y == 225) || (x == 7'd144 && y == 7'd293) || (x == 302 && y == 297) ||
		(x == 7'd569 && y == 597) || (x == 536 && y == 377) || (x == 212 && y == 281) ||
		(x == 7'd383 && y == 7'd629) || (x == 576 && y == 7'd106) || (x == 133 && y == 7'd164) ||
		(x == 7'd138 && y == 7'd461) || (x == 575 && y == 575) || (x == 292 && y == 462) ||
		(x == 131 && y == 7'd263) || (x == 223 && y == 7'd491) || (x == 7'd400 && y == 472) ||
		(x == 7'd143 && y == 7'd470) || (x == 7'd265 && y == 7'd365) || (x == 7'd432 && y == 7'd390) ||
		(x == 7'd100 && y == 593) || (x == 7'd518 && y == 7'd393) || (x == 442 && y == 273) ||
		(x == 502 && y == 216) || (x == 608 && y == 331) || (x == 7'd482 && y == 565) ||
		(x == 7'd283 && y == 172) || (x == 7'd66 && y == 634) || (x == 440 && y == 142) ||
		(x == 62 && y == 7'd303) || (x == 7'd86 && y == 7'd464) || (x == 20 && y == 7'd135) ||
		(x == 629 && y == 7'd221) || (x == 7'd119 && y == 133) || (x == 376 && y == 7'd39) ||
		(x == 147 && y == 487) || (x == 579 && y == 235) || (x == 7'd227 && y == 443) ||
		(x == 7'd238 && y == 7'd346) || (x == 7'd214 && y == 7'd345) || (x == 7'd602 && y == 273) ||
		(x == 24 && y == 7'd305) || (x == 7'd79 && y == 437) || (x == 297 && y == 364) ||
		(x == 7'd506 && y == 7'd98) || (x == 7'd621 && y == 7'd399) || (x == 482 && y == 619) ||
		(x == 521 && y == 7'd552) || (x == 625 && y == 7'd543) || (x == 224 && y == 7'd136) ||
		(x == 7'd180 && y == 7'd434) || (x == 7'd163 && y == 433) || (x == 7'd66 && y == 7'd139) ||
		(x == 7'd25 && y == 277) || (x == 516 && y == 7'd313) || (x == 7'd416 && y == 7'd402) ||
		(x == 130 && y == 7'd542) || (x == 7'd315 && y == 7'd467) || (x == 7'd468 && y == 7'd603) ||
		(x == 7'd212 && y == 249) || (x == 7'd164 && y == 7'd514) || (x == 7'd278 && y == 241) ||
		(x == 390 && y == 359) || (x == 16 && y == 7'd185) || (x == 192 && y == 7'd615) ||
		(x == 7'd572 && y == 7'd508) || (x == 460 && y == 7'd587) || (x == 294 && y == 366) ||
		(x == 7'd288 && y == 7'd466) || (x == 7'd31 && y == 168) || (x == 118 && y == 7'd524) ||
		(x == 7'd536 && y == 185) || (x == 7'd416 && y == 7'd256) || (x == 7'd215 && y == 158) ||
		(x == 558 && y == 348) || (x == 111 && y == 7'd348) || (x == 7'd385 && y == 545) ||
		(x == 502 && y == 7'd55) || (x == 638 && y == 458) || (x == 7'd272 && y == 7'd443) ||
		(x == 7'd635 && y == 27) || (x == 607 && y == 7'd59) || (x == 7'd239 && y == 349) ||
		(x == 7'd474 && y == 603) || (x == 7'd372 && y == 7'd161) || (x == 7'd389 && y == 7'd132) ||
		(x == 212 && y == 218) || (x == 7'd23 && y == 7'd264) || (x == 376 && y == 219) ||
		(x == 7'd508 && y == 318) || (x == 138 && y == 7'd408) || (x == 246 && y == 7'd582) ||
		(x == 7'd624 && y == 498) || (x == 7'd196 && y == 546) || (x == 240 && y == 7'd566) ||
		(x == 7'd348 && y == 7'd166) || (x == 636 && y == 138) || (x == 7'd343 && y == 7'd168) ||
		(x == 7'd417 && y == 7'd321) || (x == 58 && y == 7'd337) || (x == 7'd43 && y == 7'd454) ||
		(x == 211 && y == 7'd171) || (x == 344 && y == 7'd294) || (x == 7'd188 && y == 7'd270) ||
		(x == 7'd194 && y == 265) || (x == 7'd299 && y == 247) || (x == 7'd188 && y == 373) ||
		(x == 7'd69 && y == 7'd55) || (x == 7'd338 && y == 7'd568) || (x == 511 && y == 406) ||
		(x == 7'd273 && y == 7'd143) || (x == 7'd186 && y == 7'd504) || (x == 19 && y == 7'd239) ||
		(x == 224 && y == 7'd106) || (x == 7'd131 && y == 7'd379) || (x == 7'd213 && y == 311) ||
		(x == 7'd520 && y == 7'd141) || (x == 346 && y == 7'd410) || (x == 7'd8 && y == 7'd441) ||
		(x == 179 && y == 550) || (x == 7'd314 && y == 603) || (x == 7'd561 && y == 7'd354) ||
		(x == 422 && y == 633) || (x == 7'd516 && y == 7'd587) || (x == 7'd135 && y == 7'd633) ||
		(x == 7'd486 && y == 7'd5) || (x == 7'd137 && y == 7'd515) || (x == 630 && y == 327) ||
		(x == 7'd30 && y == 431) || (x == 422 && y == 7'd210) || (x == 7'd355 && y == 7'd271) ||
		(x == 250 && y == 7'd96) || (x == 159 && y == 333) || (x == 7'd322 && y == 7'd455) ||
		(x == 7'd367 && y == 19) || (x == 7'd591 && y == 7'd333) || (x == 548 && y == 188) ||
		(x == 220 && y == 625) || (x == 7'd479 && y == 504) || (x == 620 && y == 392) ||
		(x == 7'd483 && y == 7'd297) || (x == 7'd361 && y == 7'd370) || (x == 486 && y == 7'd502) ||
		(x == 232 && y == 391) || (x == 320 && y == 7'd290) || (x == 7'd388 && y == 148) ||
		(x == 7'd618 && y == 154) || (x == 609 && y == 376) || (x == 7'd622 && y == 197) ||
		(x == 7'd358 && y == 374) || (x == 448 && y == 7'd26) || (x == 63 && y == 7'd345) ||
		(x == 7'd553 && y == 439) || (x == 45 && y == 7'd125) || (x == 7'd404 && y == 7'd136) ||
		(x == 209 && y == 464) || (x == 292 && y == 7'd348) || (x == 7'd404 && y == 2) ||
		(x == 573 && y == 7'd397) || (x == 7'd495 && y == 284) || (x == 487 && y == 7'd184) ||
		(x == 349 && y == 7'd97) || (x == 7'd187 && y == 7'd525) || (x == 7'd500 && y == 7'd394) ||
		(x == 7'd295 && y == 444) || (x == 7'd437 && y == 126) || (x == 7'd92 && y == 407) ||
		(x == 7'd455 && y == 580) || (x == 363 && y == 7'd84) || (x == 7'd521 && y == 62) ||
		(x == 280 && y == 327) || (x == 7'd396 && y == 7'd244) || (x == 7'd414 && y == 7'd505) ||
		(x == 555 && y == 200) || (x == 7'd146 && y == 7'd463) || (x == 131 && y == 7'd416) ||
		(x == 312 && y == 614) || (x == 7'd222 && y == 7'd38) || (x == 7'd371 && y == 7'd389) ||
		(x == 157 && y == 7'd146) || (x == 61 && y == 7'd504) || (x == 255 && y == 7'd452) ||
		(x == 7'd5 && y == 572) || (x == 7'd286 && y == 7'd337) || (x == 231 && y == 152) ||
		(x == 7'd65 && y == 7'd305) || (x == 344 && y == 7'd212) || (x == 7'd133 && y == 7'd635) ||
		(x == 7'd122 && y == 7'd587) || (x == 571 && y == 7'd434) || (x == 7'd97 && y == 620) ||
		(x == 445 && y == 232) || (x == 178 && y == 348) || (x == 7'd446 && y == 88) ||
		(x == 7'd197 && y == 7'd270) || (x == 422 && y == 7'd438) || (x == 430 && y == 7'd383) ||
		(x == 7'd222 && y == 520) || (x == 7'd493 && y == 26) || (x == 254 && y == 7'd214) ||
		(x == 438 && y == 436) || (x == 315 && y == 573) || (x == 7'd97 && y == 547) ||
		(x == 7'd325 && y == 7'd199) || (x == 7'd599 && y == 7'd403) || (x == 7'd370 && y == 7'd453) ||
		(x == 7'd173 && y == 450) || (x == 619 && y == 7'd56) || (x == 7'd4 && y == 156) ||
		(x == 534 && y == 7'd601) || (x == 7'd609 && y == 7'd295) || (x == 485 && y == 206) ||
		(x == 333 && y == 384) || (x == 398 && y == 355) || (x == 7'd114 && y == 204) ||
		(x == 467 && y == 7'd572) || (x == 7'd506 && y == 7'd282) || (x == 7'd18 && y == 7'd448) ||
		(x == 279 && y == 7'd610) || (x == 640 && y == 533) || (x == 7'd422 && y == 584) ||
		(x == 7'd479 && y == 7'd598) || (x == 7'd365 && y == 7'd451) || (x == 7'd341 && y == 411) ||
		(x == 7'd551 && y == 7'd485) || (x == 7'd546 && y == 616) || (x == 7'd213 && y == 7'd303) ||
		(x == 547 && y == 7'd16) || (x == 257 && y == 316) || (x == 7'd358 && y == 413) ||
		(x == 7'd87 && y == 7'd386) || (x == 90 && y == 7'd239) || (x == 297 && y == 426) ||
		(x == 560 && y == 250) || (x == 536 && y == 178) || (x == 178 && y == 537) ||
		(x == 636 && y == 7'd379) || (x == 7'd64 && y == 352) || (x == 7'd273 && y == 7'd173) ||
		(x == 7'd94 && y == 7'd622) || (x == 238 && y == 501) || (x == 7'd162 && y == 7'd386) ||
		(x == 7'd381 && y == 524) || (x == 7'd188 && y == 7'd171) || (x == 7'd354 && y == 7'd327) ||
		(x == 215 && y == 510) || (x == 533 && y == 129) || (x == 7'd135 && y == 218) ||
		(x == 7'd397 && y == 7'd466) || (x == 237 && y == 7'd470) || (x == 7'd167 && y == 7'd143) ||
		(x == 281 && y == 7'd539) || (x == 460 && y == 7'd626) || (x == 7'd127 && y == 296) ||
		(x == 7'd481 && y == 7'd254) || (x == 106 && y == 99) || (x == 313 && y == 7'd532) ||
		(x == 7'd319 && y == 7'd446) || (x == 7'd398 && y == 7'd406) || (x == 457 && y == 7'd548) ||
		(x == 7'd578 && y == 124) || (x == 7'd146 && y == 37) || (x == 7'd56 && y == 454) ||
		(x == 7'd36 && y == 358) || (x == 575 && y == 377) || (x == 438 && y == 625) ||
		(x == 7'd181 && y == 563) || (x == 7'd224 && y == 508) || (x == 639 && y == 7'd596) ||
		(x == 7'd541 && y == 565) || (x == 7'd264 && y == 23) || (x == 7'd466 && y == 7'd617) ||
		(x == 65 && y == 7'd189) || (x == 7'd518 && y == 7'd433) || (x == 7'd425 && y == 7'd6) ||
		(x == 448 && y == 7'd252) || (x == 7'd332 && y == 96) || (x == 7'd48 && y == 7'd224) ||
		(x == 7'd365 && y == 7'd606) || (x == 474 && y == 559) || (x == 291 && y == 7'd535) ||
		(x == 7'd5 && y == 457) || (x == 7'd464 && y == 320) || (x == 156 && y == 7'd210) ||
		(x == 212 && y == 7'd69) || (x == 7'd403 && y == 7'd379) || (x == 501 && y == 7'd21) ||
		(x == 7'd275 && y == 7'd137) || (x == 7'd596 && y == 7'd593) || (x == 166 && y == 351) ||
		(x == 10 && y == 7'd627) || (x == 274 && y == 221) || (x == 362 && y == 7'd419) ||
		(x == 7'd291 && y == 7'd577) || (x == 7'd407 && y == 146) || (x == 7'd597 && y == 7'd598) ||
		(x == 7'd389 && y == 7'd103) || (x == 240 && y == 7'd581) || (x == 7'd198 && y == 484) ||
		(x == 234 && y == 7'd299) || (x == 7'd495 && y == 404) || (x == 7'd211 && y == 7'd283) ||
		(x == 7'd342 && y == 576) || (x == 201 && y == 567) || (x == 159 && y == 421) ||
		(x == 7'd561 && y == 7'd280) || (x == 7'd270 && y == 7'd277) || (x == 241 && y == 7'd633) ||
		(x == 7'd448 && y == 7'd47) || (x == 7'd310 && y == 7'd0) || (x == 7'd480 && y == 7'd7) ||
		(x == 574 && y == 7'd611) || (x == 596 && y == 262) || (x == 7'd131 && y == 7'd490) ||
		(x == 62 && y == 7'd426) || (x == 7'd356 && y == 7'd134) || (x == 510 && y == 478) ||
		(x == 7'd110 && y == 447) || (x == 7'd501 && y == 165) || (x == 7'd149 && y == 382) ||
		(x == 7'd523 && y == 629) || (x == 7'd46 && y == 7'd27) || (x == 7'd368 && y == 7'd16) ||
		(x == 262 && y == 483) || (x == 7'd59 && y == 7'd401) || (x == 423 && y == 7'd279) ||
		(x == 105 && y == 7'd340) || (x == 7'd383 && y == 7'd535) || (x == 7'd79 && y == 126) ||
		(x == 246 && y == 7'd556) || (x == 458 && y == 609) || (x == 417 && y == 7'd475) ||
		(x == 7'd128 && y == 455) || (x == 327 && y == 293) || (x == 7'd317 && y == 7'd44) ||
		(x == 407 && y == 449) || (x == 7'd627 && y == 7'd545) || (x == 7'd250 && y == 84) ||
		(x == 305 && y == 174) || (x == 7'd147 && y == 107) || (x == 479 && y == 7'd241) ||
		(x == 458 && y == 7'd102) || (x == 320 && y == 7'd471) || (x == 7'd20 && y == 7'd450) ||
		(x == 7'd581 && y == 7'd271) || (x == 7'd200 && y == 7'd142) || (x == 7'd593 && y == 7'd372) ||
		(x == 7'd313 && y == 129) || (x == 7'd192 && y == 517) || (x == 7'd192 && y == 7'd165) ||
		(x == 7'd24 && y == 237) || (x == 7'd133 && y == 206) || (x == 7'd8 && y == 377) ||
		(x == 7'd464 && y == 188) || (x == 7'd363 && y == 7'd152) || (x == 7'd292 && y == 7'd530) ||
		(x == 7'd207 && y == 7'd347) || (x == 422 && y == 7'd547) || (x == 7'd59 && y == 7'd345) ||
		(x == 7'd83 && y == 251) || (x == 243 && y == 7'd469) || (x == 163 && y == 164) ||
		(x == 7'd537 && y == 7'd393) || (x == 7'd369 && y == 7'd263) || (x == 312 && y == 7'd433) ||
		(x == 7'd322 && y == 7'd500) || (x == 7'd266 && y == 7'd246) || (x == 7'd534 && y == 343) ||
		(x == 67 && y == 7'd354) || (x == 7'd243 && y == 7'd58) || (x == 7'd278 && y == 464) ||
		(x == 7'd531 && y == 7'd523) || (x == 7'd393 && y == 134) || (x == 7'd615 && y == 597) ||
		(x == 7'd574 && y == 7'd55) || (x == 7'd499 && y == 7'd583) || (x == 7'd66 && y == 7'd174) ||
		(x == 7'd575 && y == 7'd596) || (x == 503 && y == 173) || (x == 489 && y == 323) ||
		(x == 635 && y == 284) || (x == 65 && y == 7'd411) || (x == 290 && y == 7'd100) ||
		(x == 341 && y == 377) || (x == 448 && y == 417) || (x == 7'd416 && y == 7'd105) ||
		(x == 439 && y == 485) || (x == 7'd145 && y == 7'd592) || (x == 633 && y == 582) ||
		(x == 7'd38 && y == 7'd146) || (x == 7'd117 && y == 7'd618) || (x == 7'd282 && y == 7'd235) ||
		(x == 7'd405 && y == 7'd538) || (x == 7'd578 && y == 9) || (x == 7'd109 && y == 248) ||
		(x == 7'd517 && y == 7'd559) || (x == 397 && y == 7'd128) || (x == 7'd178 && y == 633) ||
		(x == 133 && y == 7'd153) || (x == 7'd373 && y == 7'd393) || (x == 117 && y == 7'd313) ||
		(x == 562 && y == 7'd158) || (x == 7'd367 && y == 7'd526) || (x == 322 && y == 7'd356) ||
		(x == 7'd619 && y == 148) || (x == 7'd173 && y == 7'd361) || (x == 597 && y == 7'd96) ||
		(x == 7'd360 && y == 7'd86) || (x == 7'd547 && y == 7'd248) || (x == 218 && y == 355) ||
		(x == 7'd363 && y == 46) || (x == 7'd487 && y == 7'd330) || (x == 120 && y == 7'd418) ||
		(x == 432 && y == 393) || (x == 7'd552 && y == 631) || (x == 516 && y == 7'd76) ||
		(x == 7'd522 && y == 7'd528) || (x == 273 && y == 7'd263) || (x == 356 && y == 316) ||
		(x == 211 && y == 7'd542) || (x == 7'd387 && y == 7'd328) || (x == 7'd195 && y == 7'd293) ||
		(x == 157 && y == 7'd623) || (x == 7'd537 && y == 542) || (x == 7'd291 && y == 7'd608) ||
		(x == 166 && y == 7'd512) || (x == 7'd89 && y == 534) || (x == 7'd593 && y == 390) ||
		(x == 530 && y == 7'd80) || (x == 7'd47 && y == 7'd525) || (x == 539 && y == 7'd607) ||
		(x == 505 && y == 157) || (x == 7'd494 && y == 261) || (x == 334 && y == 7'd219) ||
		(x == 454 && y == 7'd406) || (x == 7'd316 && y == 571) || (x == 182 && y == 7'd257) ||
		(x == 7'd249 && y == 7'd232) || (x == 173 && y == 386) || (x == 7'd455 && y == 7'd133) ||
		(x == 7'd461 && y == 7'd429) || (x == 573 && y == 529) || (x == 7'd253 && y == 7'd196) ||
		(x == 565 && y == 7'd612) || (x == 300 && y == 401) || (x == 628 && y == 493) ||
		(x == 7'd321 && y == 7'd556) || (x == 226 && y == 520) || (x == 513 && y == 7'd209) ||
		(x == 216 && y == 7'd567) || (x == 7'd626 && y == 445) || (x == 461 && y == 615) ||
		(x == 227 && y == 562) || (x == 388 && y == 381) || (x == 557 && y == 427) ||
		(x == 349 && y == 599) || (x == 7'd58 && y == 7'd617) || (x == 7'd511 && y == 7'd301) ||
		(x == 297 && y == 7'd639) || (x == 7'd579 && y == 7'd498) || (x == 268 && y == 434) ||
		(x == 7'd266 && y == 7'd530) || (x == 348 && y == 410) || (x == 7'd631 && y == 38) ||
		(x == 457 && y == 7'd19) || (x == 7'd379 && y == 508) || (x == 7'd265 && y == 7'd45) ||
		(x == 228 && y == 133) || (x == 7'd579 && y == 569) || (x == 431 && y == 7'd199) ||
		(x == 7'd3 && y == 199) || (x == 7'd162 && y == 7'd451) || (x == 7'd463 && y == 341) ||
		(x == 397 && y == 622) || (x == 509 && y == 7'd575) || (x == 385 && y == 7'd149) ||
		(x == 605 && y == 7'd555) || (x == 7'd355 && y == 486) || (x == 7'd379 && y == 380) ||
		(x == 7'd522 && y == 7'd167) || (x == 7'd486 && y == 7'd199) || (x == 7'd110 && y == 539) ||
		(x == 7'd171 && y == 7'd240) || (x == 7'd110 && y == 7'd377) || (x == 7'd178 && y == 7'd589) ||
		(x == 7'd135 && y == 349) || (x == 7'd157 && y == 7'd491) || (x == 300 && y == 7'd133) ||
		(x == 359 && y == 7'd588) || (x == 388 && y == 7'd384) || (x == 7'd290 && y == 7'd215) ||
		(x == 611 && y == 579) || (x == 7'd319 && y == 7'd470) || (x == 7'd633 && y == 7'd461) ||
		(x == 193 && y == 7'd369) || (x == 7'd314 && y == 7'd259) || (x == 7'd626 && y == 7'd165) ||
		(x == 517 && y == 467) || (x == 7'd597 && y == 7'd583) || (x == 7'd21 && y == 7'd288) ||
		(x == 195 && y == 456) || (x == 7'd151 && y == 230) || (x == 7'd510 && y == 7'd210) ||
		(x == 7'd408 && y == 7'd390) || (x == 7'd297 && y == 7'd524) || (x == 7'd342 && y == 334) ||
		(x == 515 && y == 443) || (x == 7'd332 && y == 7'd33) || (x == 379 && y == 7'd179) ||
		(x == 7'd110 && y == 7'd5) || (x == 227 && y == 410) || (x == 436 && y == 7'd507) ||
		(x == 7'd238 && y == 7'd258) || (x == 470 && y == 7'd598) || (x == 221 && y == 252) ||
		(x == 297 && y == 7'd47) || (x == 330 && y == 436) || (x == 7'd605 && y == 605) ||
		(x == 7'd604 && y == 7'd382) || (x == 220 && y == 7'd45) || (x == 7'd493 && y == 7'd598) ||
		(x == 7'd246 && y == 7'd365) || (x == 412 && y == 170) || (x == 7'd425 && y == 7'd387) ||
		(x == 7'd572 && y == 136) || (x == 7'd306 && y == 7'd617) || (x == 7'd3 && y == 616) ||
		(x == 7'd354 && y == 140) || (x == 7'd461 && y == 239) || (x == 7'd448 && y == 7'd343) ||
		(x == 7'd113 && y == 7'd368) || (x == 229 && y == 7'd350) || (x == 7'd407 && y == 181) ||
		(x == 7'd57 && y == 259) || (x == 183 && y == 7'd282) || (x == 7'd593 && y == 105) ||
		(x == 311 && y == 7'd375) || (x == 7'd484 && y == 7'd618) || (x == 519 && y == 7'd197) ||
		(x == 7'd486 && y == 227) || (x == 7'd477 && y == 461) || (x == 457 && y == 546) ||
		(x == 321 && y == 7'd179) || (x == 454 && y == 7'd10) || (x == 166 && y == 7'd99) ||
		(x == 7'd245 && y == 7'd237) || (x == 7'd221 && y == 357) || (x == 515 && y == 7'd569) ||
		(x == 206 && y == 7'd423) || (x == 7'd185 && y == 7'd341) || (x == 7'd368 && y == 38) ||
		(x == 474 && y == 502) || (x == 216 && y == 582) || (x == 489 && y == 7'd120) ||
		(x == 7'd615 && y == 7'd259) || (x == 513 && y == 7'd406) || (x == 7'd597 && y == 430) ||
		(x == 7'd246 && y == 7'd597) || (x == 431 && y == 609) || (x == 346 && y == 7'd26) ||
		(x == 7'd534 && y == 7'd264) || (x == 7'd16 && y == 7'd567) || (x == 55 && y == 7'd453) ||
		(x == 7'd611 && y == 518) || (x == 7'd613 && y == 7'd253) || (x == 7'd66 && y == 260) ||
		(x == 544 && y == 7'd157) || (x == 7'd550 && y == 7'd355) || (x == 7'd572 && y == 7'd261) ||
		(x == 7'd373 && y == 248) || (x == 7'd336 && y == 578) || (x == 7'd404 && y == 3) ||
		(x == 7'd170 && y == 603) || (x == 408 && y == 7'd372) || (x == 7'd624 && y == 283) ||
		(x == 197 && y == 193) || (x == 7'd482 && y == 7'd620) || (x == 7'd529 && y == 7'd630) ||
		(x == 7'd574 && y == 7'd194) || (x == 542 && y == 7'd260) || (x == 7'd322 && y == 7'd370) ||
		(x == 472 && y == 201) || (x == 7'd524 && y == 7'd462) || (x == 273 && y == 341) ||
		(x == 7'd65 && y == 7'd298) || (x == 361 && y == 324) || (x == 7'd539 && y == 7'd3) ||
		(x == 447 && y == 7'd170) || (x == 256 && y == 7'd185) || (x == 7'd572 && y == 7'd258) ||
		(x == 519 && y == 636) || (x == 7'd93 && y == 155) || (x == 7'd290 && y == 419) ||
		(x == 485 && y == 479) || (x == 7'd225 && y == 7'd305) || (x == 7'd482 && y == 7'd8) ||
		(x == 7'd344 && y == 7'd261) || (x == 7'd368 && y == 474) || (x == 373 && y == 436) ||
		(x == 17 && y == 7'd450) || (x == 609 && y == 274) || (x == 508 && y == 7'd345) ||
		(x == 7'd293 && y == 7'd627) || (x == 7'd366 && y == 7'd497) || (x == 7'd321 && y == 498) ||
		(x == 583 && y == 545) || (x == 301 && y == 7'd271) || (x == 7'd560 && y == 191) ||
		(x == 364 && y == 7'd274) || (x == 148 && y == 614) || (x == 7'd159 && y == 313) ||
		(x == 453 && y == 406) || (x == 552 && y == 530) || (x == 7'd385 && y == 608) ||
		(x == 635 && y == 7'd322) || (x == 239 && y == 472) || (x == 7'd197 && y == 7'd459) ||
		(x == 7'd36 && y == 140) || (x == 198 && y == 250) || (x == 420 && y == 7'd541) ||
		(x == 7'd619 && y == 403) || (x == 250 && y == 143) || (x == 7'd453 && y == 7'd520) ||
		(x == 7'd529 && y == 7'd556) || (x == 7'd620 && y == 7'd297) || (x == 83 && y == 7'd556) ||
		(x == 7'd601 && y == 7'd8) || (x == 306 && y == 142) || (x == 7'd227 && y == 7'd436) ||
		(x == 7'd147 && y == 7'd568) || (x == 615 && y == 7'd241) || (x == 7'd400 && y == 7'd237) ||
		(x == 7'd81 && y == 115) || (x == 501 && y == 7'd95) || (x == 7'd190 && y == 7'd582) ||
		(x == 7'd193 && y == 7'd235) || (x == 7'd16 && y == 7'd240) || (x == 7'd329 && y == 7'd462) ||
		(x == 384 && y == 7'd612) || (x == 7'd142 && y == 7'd65) || (x == 7'd103 && y == 393) ||
		(x == 7'd347 && y == 7'd38) || (x == 171 && y == 569) || (x == 7'd393 && y == 465) ||
		(x == 7'd500 && y == 7'd586) || (x == 201 && y == 7'd163) || (x == 7'd34 && y == 636) ||
		(x == 176 && y == 7'd382) || (x == 245 && y == 7'd189) || (x == 7'd621 && y == 7'd578) ||
		(x == 427 && y == 7'd592) || (x == 7'd235 && y == 7'd375) || (x == 7'd271 && y == 7'd369) ||
		(x == 7'd618 && y == 7'd455) || (x == 7'd398 && y == 7'd628) || (x == 7'd588 && y == 609) ||
		(x == 166 && y == 239) || (x == 623 && y == 546) || (x == 7'd525 && y == 182) ||
		(x == 7'd365 && y == 294) || (x == 580 && y == 378) || (x == 7'd449 && y == 63) ||
		(x == 7'd68 && y == 7'd208) || (x == 7'd230 && y == 7'd237) || (x == 548 && y == 363) ||
		(x == 7'd423 && y == 472) || (x == 363 && y == 7'd580) || (x == 7'd132 && y == 308) ||
		(x == 7'd153 && y == 399) || (x == 260 && y == 156) || (x == 7'd540 && y == 7'd107) ||
		(x == 577 && y == 7'd416) || (x == 7'd484 && y == 378) || (x == 7'd571 && y == 7'd87) ||
		(x == 7'd151 && y == 556) || (x == 7'd238 && y == 495) || (x == 7'd151 && y == 51) ||
		(x == 7'd470 && y == 7'd120) || (x == 7'd380 && y == 184) || (x == 7'd205 && y == 498) ||
		(x == 464 && y == 382) || (x == 190 && y == 7'd177) || (x == 197 && y == 7'd496) ||
		(x == 616 && y == 435) || (x == 324 && y == 616) || (x == 7'd218 && y == 7'd419) ||
		(x == 7'd636 && y == 7'd271) || (x == 587 && y == 7'd25) || (x == 7'd536 && y == 7'd126) ||
		(x == 7'd224 && y == 7'd424) || (x == 593 && y == 496) || (x == 7'd507 && y == 7'd631) ||
		(x == 318 && y == 418) || (x == 7'd453 && y == 7'd510) || (x == 213 && y == 7'd596) ||
		(x == 7'd377 && y == 571) || (x == 7'd118 && y == 7'd327) || (x == 7'd253 && y == 7'd619) ||
		(x == 602 && y == 7'd49) || (x == 527 && y == 462) || (x == 182 && y == 452) ||
		(x == 7'd528 && y == 23) || (x == 322 && y == 7'd90) || (x == 7'd534 && y == 7'd76) ||
		(x == 361 && y == 387) || (x == 7'd368 && y == 32) || (x == 439 && y == 504) ||
		(x == 419 && y == 560) || (x == 7'd622 && y == 406) || (x == 347 && y == 355) ||
		(x == 7'd171 && y == 582) || (x == 175 && y == 7'd55) || (x == 7'd590 && y == 7'd512) ||
		(x == 7'd207 && y == 212) || (x == 7'd338 && y == 202) || (x == 120 && y == 7'd413) ||
		(x == 7'd154 && y == 184) || (x == 319 && y == 434) || (x == 7'd618 && y == 7'd153) ||
		(x == 401 && y == 181) || (x == 167 && y == 7'd316) || (x == 345 && y == 7'd321) ||
		(x == 7'd390 && y == 7'd302) || (x == 232 && y == 7'd569) || (x == 434 && y == 7'd80) ||
		(x == 7'd74 && y == 7'd404) || (x == 7'd593 && y == 293) || (x == 240 && y == 161) ||
		(x == 7'd498 && y == 7'd382) || (x == 7'd413 && y == 7'd588) || (x == 7'd159 && y == 7'd467) ||
		(x == 7'd114 && y == 7'd132) || (x == 7'd303 && y == 465) || (x == 7'd20 && y == 631) ||
		(x == 89 && y == 7'd528) || (x == 7'd611 && y == 7'd487) || (x == 424 && y == 183) ||
		(x == 7'd471 && y == 202) || (x == 7'd198 && y == 7'd590) || (x == 7'd143 && y == 37) ||
		(x == 465 && y == 7'd193) || (x == 7'd475 && y == 7'd390) || (x == 192 && y == 216) ||
		(x == 460 && y == 441) || (x == 103 && y == 125) || (x == 7'd52 && y == 208) ||
		(x == 243 && y == 7'd487) || (x == 599 && y == 7'd399) || (x == 306 && y == 540) ||
		(x == 239 && y == 7'd314) || (x == 7'd581 && y == 216) || (x == 7'd496 && y == 7'd391) ||
		(x == 405 && y == 196) || (x == 7'd627 && y == 7'd421) || (x == 7'd293 && y == 613) ||
		(x == 436 && y == 577) || (x == 7'd238 && y == 499) || (x == 606 && y == 370) ||
		(x == 7'd622 && y == 268) || (x == 574 && y == 494) || (x == 231 && y == 7'd563) ||
		(x == 301 && y == 7'd441) || (x == 7'd306 && y == 7'd401) || (x == 7'd635 && y == 7'd123) ||
		(x == 7'd420 && y == 7'd472) || (x == 7'd247 && y == 7'd399) || (x == 131 && y == 7'd273) ||
		(x == 7'd81 && y == 7'd248) || (x == 153 && y == 7'd579) || (x == 7'd219 && y == 157) ||
		(x == 13 && y == 7'd80) || (x == 7'd124 && y == 7'd564) || (x == 569 && y == 7'd78) ||
		(x == 278 && y == 7'd291) || (x == 317 && y == 544) || (x == 7'd41 && y == 7'd567) ||
		(x == 7'd192 && y == 436) || (x == 238 && y == 519) || (x == 514 && y == 7'd553) ||
		(x == 149 && y == 639) || (x == 576 && y == 393) || (x == 7'd365 && y == 7'd246) ||
		(x == 7'd243 && y == 525) || (x == 438 && y == 475) || (x == 7'd179 && y == 7'd486) ||
		(x == 495 && y == 7'd84) || (x == 633 && y == 7'd78) || (x == 278 && y == 7'd371) ||
		(x == 7'd254 && y == 7'd276) || (x == 7'd393 && y == 7'd117) || (x == 342 && y == 7'd590) ||
		(x == 7'd627 && y == 7'd348) || (x == 521 && y == 7'd426) || (x == 67 && y == 7'd591) ||
		(x == 462 && y == 7'd133) || (x == 480 && y == 357) || (x == 7'd369 && y == 7'd313) ||
		(x == 7'd318 && y == 7'd631) || (x == 198 && y == 605) || (x == 7'd321 && y == 289) ||
		(x == 320 && y == 7'd423) || (x == 476 && y == 7'd109) || (x == 272 && y == 7'd591) ||
		(x == 3 && y == 7'd432) || (x == 7'd145 && y == 7'd596) || (x == 7'd384 && y == 354) ||
		(x == 7'd380 && y == 449) || (x == 478 && y == 7'd422) || (x == 7'd429 && y == 436) ||
		(x == 7'd311 && y == 7'd468) || (x == 7'd46 && y == 171) || (x == 7'd203 && y == 300) ||
		(x == 7'd570 && y == 83) || (x == 265 && y == 7'd187) || (x == 7'd493 && y == 7'd144) ||
		(x == 7'd190 && y == 7'd400) || (x == 7'd339 && y == 561) || (x == 524 && y == 7'd256) ||
		(x == 7'd581 && y == 569) || (x == 7'd20 && y == 118) || (x == 7'd277 && y == 502) ||
		(x == 343 && y == 191) || (x == 274 && y == 7'd17) || (x == 7'd536 && y == 382) ||
		(x == 559 && y == 333) || (x == 376 && y == 314) || (x == 89 && y == 7'd414) ||
		(x == 7'd518 && y == 1) || (x == 7'd327 && y == 416) || (x == 7'd495 && y == 7'd219) ||
		(x == 88 && y == 7'd391) || (x == 7'd405 && y == 7'd559) || (x == 7'd358 && y == 7'd510) ||
		(x == 59 && y == 7'd380) || (x == 224 && y == 229) || (x == 332 && y == 562) ||
		(x == 7'd635 && y == 7'd308) || (x == 576 && y == 525) || (x == 7'd467 && y == 7'd180) ||
		(x == 7'd449 && y == 7'd432) || (x == 279 && y == 366) || (x == 144 && y == 7'd117) ||
		(x == 223 && y == 7'd312) || (x == 7'd309 && y == 20) || (x == 292 && y == 331) ||
		(x == 7'd382 && y == 415) || (x == 7'd338 && y == 457) || (x == 7'd255 && y == 463) ||
		(x == 635 && y == 530) || (x == 7'd134 && y == 7'd517) || (x == 7'd39 && y == 7'd233) ||
		(x == 165 && y == 224) || (x == 321 && y == 7'd253) || (x == 7'd581 && y == 7'd352) ||
		(x == 7'd298 && y == 7'd268) || (x == 7'd481 && y == 194) || (x == 7'd553 && y == 7'd375) ||
		(x == 7'd505 && y == 108) || (x == 7'd196 && y == 7'd516) || (x == 7'd187 && y == 145) ||
		(x == 103 && y == 7'd4) || (x == 7'd624 && y == 291) || (x == 406 && y == 182) ||
		(x == 7'd144 && y == 7'd316) || (x == 7'd466 && y == 125) || (x == 7'd399 && y == 7'd426) ||
		(x == 347 && y == 7'd96) || (x == 340 && y == 7'd212) || (x == 7'd343 && y == 485) ||
		(x == 199 && y == 7'd37) || (x == 103 && y == 7'd431) || (x == 7'd529 && y == 7'd565) ||
		(x == 70 && y == 7'd587) || (x == 7'd228 && y == 7'd363) || (x == 596 && y == 7'd130) ||
		(x == 7'd626 && y == 454) || (x == 7'd140 && y == 319) || (x == 163 && y == 185) ||
		(x == 141 && y == 7'd153) || (x == 472 && y == 611) || (x == 600 && y == 7'd576) ||
		(x == 7'd504 && y == 7'd397) || (x == 7'd125 && y == 7'd413) || (x == 36 && y == 7'd631) ||
		(x == 7'd375 && y == 507) || (x == 298 && y == 310) || (x == 7'd383 && y == 287) ||
		(x == 7'd74 && y == 615) || (x == 7'd626 && y == 7'd216) || (x == 7'd500 && y == 7'd98) ||
		(x == 7'd620 && y == 7'd556) || (x == 488 && y == 7'd116) || (x == 639 && y == 231) ||
		(x == 7'd505 && y == 418) || (x == 7'd103 && y == 476) || (x == 192 && y == 418) ||
		(x == 7'd288 && y == 7'd299) || (x == 7'd588 && y == 84) || (x == 341 && y == 7'd633) ||
		(x == 7'd344 && y == 134) || (x == 7'd118 && y == 7'd87) || (x == 630 && y == 7'd253) ||
		(x == 595 && y == 7'd288) || (x == 612 && y == 313) || (x == 7'd225 && y == 624) ||
		(x == 7'd579 && y == 7'd499) || (x == 7'd264 && y == 1) || (x == 115 && y == 7'd324) ||
		(x == 7'd447 && y == 7'd348) || (x == 429 && y == 7'd110) || (x == 7'd486 && y == 7'd552) ||
		(x == 7'd524 && y == 157) || (x == 276 && y == 7'd194) || (x == 245 && y == 573) ||
		(x == 324 && y == 7'd14) || (x == 21 && y == 7'd11) || (x == 561 && y == 501) ||
		(x == 7'd445 && y == 7'd261) || (x == 7'd54 && y == 7'd105) || (x == 7'd251 && y == 7'd154) ||
		(x == 7'd610 && y == 7'd618) || (x == 318 && y == 7'd150) || (x == 580 && y == 163) ||
		(x == 68 && y == 7'd494) || (x == 249 && y == 7'd113) || (x == 7'd485 && y == 342) ||
		(x == 498 && y == 7'd564) || (x == 593 && y == 7'd446) || (x == 305 && y == 7'd286) ||
		(x == 353 && y == 540) || (x == 114 && y == 7'd201) || (x == 7'd472 && y == 404) ||
		(x == 267 && y == 7'd57) || (x == 7'd98 && y == 7'd550) || (x == 7'd138 && y == 7'd420) ||
		(x == 499 && y == 339) || (x == 7'd55 && y == 494) || (x == 621 && y == 141) ||
		(x == 7'd64 && y == 532) || (x == 556 && y == 7'd356) || (x == 7'd309 && y == 7'd401) ||
		(x == 130 && y == 629) || (x == 7'd135 && y == 7'd536) || (x == 7'd96 && y == 162) ||
		(x == 186 && y == 7'd117) || (x == 7'd317 && y == 7'd340) || (x == 7'd49 && y == 187) ||
		(x == 7'd261 && y == 317) || (x == 434 && y == 7'd89) || (x == 460 && y == 251) ||
		(x == 311 && y == 7'd527) || (x == 7'd150 && y == 7'd178) || (x == 159 && y == 7'd404) ||
		(x == 591 && y == 406) || (x == 7'd253 && y == 7'd227) || (x == 7'd596 && y == 347) ||
		(x == 428 && y == 7'd579) || (x == 565 && y == 7'd361) || (x == 7'd366 && y == 547) ||
		(x == 7'd116 && y == 7'd524) || (x == 7'd521 && y == 7'd494) || (x == 7'd111 && y == 7'd269) ||
		(x == 321 && y == 7'd447) || (x == 575 && y == 227) || (x == 7'd625 && y == 7'd436) ||
		(x == 413 && y == 592) || (x == 7'd205 && y == 7'd171) || (x == 7'd354 && y == 154) ||
		(x == 7'd206 && y == 7'd233) || (x == 7'd343 && y == 591) || (x == 7'd155 && y == 519) ||
		(x == 7'd254 && y == 7'd149) || (x == 112 && y == 7'd143) || (x == 62 && y == 7'd390) ||
		(x == 7'd92 && y == 445) || (x == 7'd223 && y == 546) || (x == 344 && y == 7'd27) ||
		(x == 490 && y == 456) || (x == 7'd204 && y == 7'd16) || (x == 192 && y == 590) ||
		(x == 383 && y == 7'd614) || (x == 7'd234 && y == 7'd513) || (x == 529 && y == 7'd550) ||
		(x == 7'd262 && y == 7'd130) || (x == 7'd318 && y == 7'd413) || (x == 427 && y == 411) ||
		(x == 7'd244 && y == 345) || (x == 7'd626 && y == 7'd290) || (x == 595 && y == 200) ||
		(x == 7'd539 && y == 7'd565) || (x == 388 && y == 7'd579) || (x == 314 && y == 224) ||
		(x == 433 && y == 7'd243) || (x == 7'd454 && y == 591) || (x == 145 && y == 160) ||
		(x == 487 && y == 7'd545) || (x == 7'd344 && y == 7'd18) || (x == 580 && y == 276) ||
		(x == 166 && y == 477) || (x == 335 && y == 7'd380) || (x == 7'd634 && y == 7'd209) ||
		(x == 181 && y == 193) || (x == 7'd382 && y == 7'd357) || (x == 7'd325 && y == 7'd569) ||
		(x == 7'd295 && y == 305) || (x == 389 && y == 7'd547) || (x == 7'd615 && y == 331) ||
		(x == 190 && y == 596) || (x == 574 && y == 7'd552) || (x == 7'd358 && y == 431) ||
		(x == 7'd554 && y == 7'd252) || (x == 307 && y == 186) || (x == 245 && y == 7'd255) ||
		(x == 7'd368 && y == 252) || (x == 244 && y == 7'd246) || (x == 323 && y == 267) ||
		(x == 7'd190 && y == 7'd397) || (x == 616 && y == 456) || (x == 191 && y == 7'd377) ||
		(x == 7'd260 && y == 25) || (x == 7'd404 && y == 7'd517) || (x == 7'd135 && y == 7'd375) ||
		(x == 7'd594 && y == 7'd240) || (x == 15 && y == 7'd599) || (x == 7'd217 && y == 7'd424) ||
		(x == 416 && y == 376) || (x == 640 && y == 7'd440) || (x == 7'd96 && y == 531) ||
		(x == 7'd73 && y == 351) || (x == 7'd277 && y == 307) || (x == 7'd547 && y == 381) ||
		(x == 562 && y == 7'd193) || (x == 615 && y == 559) || (x == 283 && y == 7'd346) ||
		(x == 7'd327 && y == 7'd330) || (x == 253 && y == 548) || (x == 7'd382 && y == 53) ||
		(x == 7'd487 && y == 7'd468) || (x == 7'd574 && y == 7'd514) || (x == 7'd33 && y == 310) ||
		(x == 493 && y == 7'd296) || (x == 7'd410 && y == 7'd515) || (x == 7'd375 && y == 483) ||
		(x == 7'd542 && y == 7'd339) || (x == 7'd145 && y == 7'd448) || (x == 7'd349 && y == 7'd236) ||
		(x == 400 && y == 7'd257) || (x == 407 && y == 7'd412) || (x == 7'd342 && y == 153) ||
		(x == 7'd406 && y == 7'd409) || (x == 205 && y == 7'd278) || (x == 309 && y == 7'd412) ||
		(x == 7'd248 && y == 7'd549) || (x == 482 && y == 7'd473) || (x == 7'd111 && y == 88) ||
		(x == 490 && y == 314) || (x == 7'd582 && y == 7'd156) || (x == 393 && y == 7'd259) ||
		(x == 7'd262 && y == 7'd30) || (x == 7'd376 && y == 7'd236) || (x == 275 && y == 7'd548) ||
		(x == 7'd41 && y == 341) || (x == 507 && y == 455) || (x == 7'd530 && y == 400) ||
		(x == 268 && y == 398) || (x == 7'd196 && y == 7'd184) || (x == 299 && y == 7'd11) ||
		(x == 7'd554 && y == 7'd408) || (x == 7'd490 && y == 7'd258) || (x == 7'd605 && y == 7'd539) ||
		(x == 7'd326 && y == 421) || (x == 7'd199 && y == 36) || (x == 7'd150 && y == 7'd538) ||
		(x == 55 && y == 7'd467) || (x == 7'd344 && y == 7'd283) || (x == 7'd571 && y == 7'd28) ||
		(x == 596 && y == 366) || (x == 483 && y == 7'd358) || (x == 290 && y == 143) ||
		(x == 7'd318 && y == 622) || (x == 7'd461 && y == 7'd339) || (x == 7'd368 && y == 234) ||
		(x == 151 && y == 7'd188) || (x == 7'd290 && y == 577) || (x == 467 && y == 7'd284) ||
		(x == 355 && y == 7'd141) || (x == 11 && y == 7'd315) || (x == 7'd122 && y == 561) ||
		(x == 7'd293 && y == 7'd389) || (x == 304 && y == 7'd225) || (x == 7'd342 && y == 7'd260) ||
		(x == 546 && y == 620) || (x == 319 && y == 7'd321) || (x == 7'd71 && y == 7'd332) ||
		(x == 7'd630 && y == 7'd364) || (x == 452 && y == 370) || (x == 7'd377 && y == 7'd515) ||
		(x == 7'd138 && y == 81) || (x == 7'd401 && y == 7'd406) || (x == 516 && y == 7'd196) ||
		(x == 7'd28 && y == 7'd436) || (x == 7'd22 && y == 7) || (x == 7'd136 && y == 7'd256) ||
		(x == 7'd241 && y == 626) || (x == 7'd320 && y == 7'd188) || (x == 7'd197 && y == 7'd338) ||
		(x == 126 && y == 7'd155) || (x == 7'd537 && y == 532) || (x == 7'd621 && y == 323) ||
		(x == 7'd190 && y == 7'd341) || (x == 7'd412 && y == 7'd350) || (x == 625 && y == 7'd502) ||
		(x == 7'd630 && y == 7'd36) || (x == 232 && y == 488) || (x == 7'd189 && y == 7'd15) ||
		(x == 495 && y == 613) || (x == 174 && y == 7'd431) || (x == 7'd393 && y == 7'd524) ||
		(x == 7'd3 && y == 7'd482) || (x == 7'd247 && y == 321) || (x == 492 && y == 7'd569) ||
		(x == 7'd597 && y == 7'd506) || (x == 7'd121 && y == 7'd414) || (x == 407 && y == 368) ||
		(x == 7'd550 && y == 276) || (x == 7'd16 && y == 7'd294) || (x == 393 && y == 583) ||
		(x == 7'd115 && y == 7'd636) || (x == 7'd625 && y == 7'd439) || (x == 7'd518 && y == 430) ||
		(x == 7'd550 && y == 7'd503) || (x == 90 && y == 7'd509) || (x == 473 && y == 7'd481) ||
		(x == 197 && y == 204) || (x == 292 && y == 7'd585) || (x == 423 && y == 296) ||
		(x == 256 && y == 498) || (x == 7'd492 && y == 272) || (x == 7'd212 && y == 414) ||
		(x == 395 && y == 602) || (x == 7'd313 && y == 7'd233) || (x == 229 && y == 345) ||
		(x == 7'd108 && y == 7'd296) || (x == 154 && y == 7'd562) || (x == 7'd603 && y == 7'd506) ||
		(x == 41 && y == 7'd49) || (x == 521 && y == 433) || (x == 315 && y == 7'd487) ||
		(x == 28 && y == 7'd259) || (x == 7'd280 && y == 414) || (x == 7'd272 && y == 7'd289) ||
		(x == 7'd367 && y == 7'd41) || (x == 358 && y == 568) || (x == 7'd15 && y == 455) ||
		(x == 331 && y == 7'd348) || (x == 7'd174 && y == 538) || (x == 7'd388 && y == 614) ||
		(x == 210 && y == 7'd491) || (x == 7'd132 && y == 7'd520) || (x == 203 && y == 7'd476) ||
		(x == 7'd143 && y == 386) || (x == 314 && y == 7'd433) || (x == 7'd467 && y == 7'd379) ||
		(x == 7'd283 && y == 413) || (x == 393 && y == 7'd129) || (x == 7'd245 && y == 123) ||
		(x == 580 && y == 7'd277) || (x == 7'd619 && y == 120) || (x == 7'd112 && y == 494) ||
		(x == 7'd398 && y == 7'd169) || (x == 7'd529 && y == 358) || (x == 500 && y == 354) ||
		(x == 541 && y == 7'd42) || (x == 7'd623 && y == 191) || (x == 7'd251 && y == 7'd263) ||
		(x == 7'd27 && y == 371) || (x == 7'd68 && y == 611) || (x == 186 && y == 305) ||
		(x == 529 && y == 432) || (x == 612 && y == 638) || (x == 7'd533 && y == 7'd633) ||
		(x == 7'd26 && y == 521) || (x == 7'd389 && y == 7'd304) || (x == 7'd241 && y == 7'd631) ||
		(x == 7'd242 && y == 7'd87) || (x == 7'd478 && y == 7'd254) || (x == 364 && y == 575) ||
		(x == 138 && y == 463) || (x == 637 && y == 267) || (x == 7'd564 && y == 40) ||
		(x == 418 && y == 313) || (x == 416 && y == 7'd298) || (x == 416 && y == 578) ||
		(x == 7'd305 && y == 208) || (x == 628 && y == 400) || (x == 493 && y == 556) ||
		(x == 7'd303 && y == 396) || (x == 396 && y == 582) || (x == 7'd575 && y == 7'd631) ||
		(x == 7'd548 && y == 398) || (x == 370 && y == 328) || (x == 7'd462 && y == 7'd254) ||
		(x == 527 && y == 608) || (x == 7'd167 && y == 7'd317) || (x == 512 && y == 7'd433) ||
		(x == 370 && y == 7'd446) || (x == 7'd467 && y == 7'd443) || (x == 7'd33 && y == 143) ||
		(x == 149 && y == 136) || (x == 443 && y == 7'd154) || (x == 7'd240 && y == 7'd367) ||
		(x == 7'd410 && y == 7'd537) || (x == 7'd467 && y == 7'd582) || (x == 7'd564 && y == 543) ||
		(x == 7'd253 && y == 7'd556) || (x == 7'd596 && y == 7'd387) || (x == 7'd193 && y == 7'd633) ||
		(x == 7'd130 && y == 7'd634) || (x == 275 && y == 255) || (x == 7'd445 && y == 7'd351) ||
		(x == 327 && y == 440) || (x == 619 && y == 575) || (x == 7'd552 && y == 10) ||
		(x == 7'd523 && y == 7'd43) || (x == 335 && y == 7'd190) || (x == 7'd448 && y == 7'd557) ||
		(x == 192 && y == 7'd481) || (x == 202 && y == 7'd400) || (x == 7'd246 && y == 60) ||
		(x == 7'd140 && y == 7'd42) || (x == 7'd396 && y == 7'd214) || (x == 463 && y == 7'd115) ||
		(x == 7'd404 && y == 7'd492) || (x == 7'd547 && y == 7'd631) || (x == 7'd236 && y == 84) ||
		(x == 7'd605 && y == 628) || (x == 467 && y == 7'd604) || (x == 7'd488 && y == 7'd614) ||
		(x == 7'd312 && y == 317) || (x == 7'd467 && y == 7'd173) || (x == 426 && y == 7'd305) ||
		(x == 111 && y == 7'd298) || (x == 7'd342 && y == 7'd354) || (x == 366 && y == 430) ||
		(x == 120 && y == 7'd395) || (x == 7'd630 && y == 7'd481) || (x == 7'd87 && y == 7'd260) ||
		(x == 7'd576 && y == 7'd262) || (x == 292 && y == 615) || (x == 260 && y == 7'd126) ||
		(x == 7'd14 && y == 7'd213) || (x == 7'd460 && y == 7'd181) || (x == 7'd63 && y == 277) ||
		(x == 158 && y == 7'd425) || (x == 478 && y == 505) || (x == 555 && y == 7'd308) ||
		(x == 7'd513 && y == 236) || (x == 7'd479 && y == 7'd144) || (x == 7'd511 && y == 7'd309) ||
		(x == 370 && y == 197) || (x == 7'd302 && y == 474) || (x == 7'd210 && y == 7'd58) ||
		(x == 7'd466 && y == 7'd578) || (x == 7'd385 && y == 193) || (x == 448 && y == 362) ||
		(x == 7'd584 && y == 7'd390) || (x == 7'd154 && y == 307) || (x == 150 && y == 153) ||
		(x == 7'd137 && y == 342) || (x == 277 && y == 543) || (x == 190 && y == 7'd439) ||
		(x == 7'd214 && y == 7'd295) || (x == 7'd359 && y == 7'd146) || (x == 334 && y == 7'd612) ||
		(x == 622 && y == 309) || (x == 592 && y == 463) || (x == 7'd380 && y == 7'd78) ||
		(x == 7'd619 && y == 7'd611) || (x == 185 && y == 213) || (x == 7'd556 && y == 7'd519) ||
		(x == 7'd624 && y == 228) || (x == 391 && y == 7'd340) || (x == 7'd189 && y == 273) ||
		(x == 7'd529 && y == 7'd111) || (x == 18 && y == 7'd278) || (x == 190 && y == 638) ||
		(x == 7'd253 && y == 7'd233) || (x == 271 && y == 7'd240) || (x == 7'd486 && y == 302) ||
		(x == 291 && y == 7'd305) || (x == 7'd374 && y == 56) || (x == 7'd405 && y == 7'd521) ||
		(x == 7'd508 && y == 387) || (x == 76 && y == 7'd301) || (x == 124 && y == 7'd614) ||
		(x == 191 && y == 343) || (x == 474 && y == 7'd51) || (x == 294 && y == 7'd387) ||
		(x == 7'd238 && y == 469) || (x == 634 && y == 7'd511) || (x == 493 && y == 7'd537) ||
		(x == 7'd495 && y == 7'd39) || (x == 7'd443 && y == 7'd142) || (x == 212 && y == 418) ||
		(x == 7'd360 && y == 551) || (x == 7'd445 && y == 502) || (x == 212 && y == 7'd378) ||
		(x == 7'd79 && y == 636) || (x == 7'd637 && y == 7'd231) || (x == 568 && y == 7'd439) ||
		(x == 15 && y == 7'd143) || (x == 613 && y == 514) || (x == 7'd547 && y == 7'd489) ||
		(x == 412 && y == 302) || (x == 7'd304 && y == 276) || (x == 566 && y == 7'd458) ||
		(x == 7'd191 && y == 7'd471) || (x == 7'd344 && y == 193) || (x == 334 && y == 213) ||
		(x == 275 && y == 262) || (x == 375 && y == 218) || (x == 7'd616 && y == 182) ||
		(x == 628 && y == 483) || (x == 7'd223 && y == 7'd327) || (x == 7'd351 && y == 327) ||
		(x == 7'd452 && y == 7'd267) || (x == 245 && y == 7'd371) || (x == 137 && y == 156) ||
		(x == 7'd555 && y == 7'd39) || (x == 7'd157 && y == 7'd528) || (x == 456 && y == 7'd216) ||
		(x == 7'd462 && y == 421) || (x == 7'd467 && y == 7'd184) || (x == 7'd275 && y == 266) ||
		(x == 7'd542 && y == 7'd156) || (x == 7'd628 && y == 7'd369) || (x == 247 && y == 405) ||
		(x == 69 && y == 7'd206) || (x == 372 && y == 427) || (x == 7'd543 && y == 44) ||
		(x == 7'd417 && y == 7'd217) || (x == 7'd600 && y == 7'd241) || (x == 7'd424 && y == 7'd238) ||
		(x == 218 && y == 563) || (x == 7'd368 && y == 338) || (x == 7'd602 && y == 7'd290) ||
		(x == 183 && y == 543) || (x == 7'd209 && y == 342) || (x == 7'd360 && y == 115) ||
		(x == 370 && y == 207) || (x == 426 && y == 613) || (x == 307 && y == 7'd625) ||
		(x == 543 && y == 7'd65) || (x == 320 && y == 506) || (x == 455 && y == 7'd563) ||
		(x == 489 && y == 389) || (x == 638 && y == 7'd469) || (x == 265 && y == 7'd526) ||
		(x == 7'd402 && y == 478) || (x == 302 && y == 7'd73) || (x == 140 && y == 568) ||
		(x == 160 && y == 7'd21) || (x == 191 && y == 7'd54) || (x == 7'd293 && y == 7'd13) ||
		(x == 237 && y == 7'd134) || (x == 465 && y == 7'd534) || (x == 503 && y == 523) ||
		(x == 7'd189 && y == 7'd447) || (x == 414 && y == 7'd539) || (x == 7'd16 && y == 7'd596) ||
		(x == 598 && y == 7'd341) || (x == 7'd231 && y == 609) || (x == 7'd333 && y == 7'd207) ||
		(x == 145 && y == 336) || (x == 7'd109 && y == 7'd631) || (x == 460 && y == 637) ||
		(x == 84 && y == 7'd105) || (x == 168 && y == 520) || (x == 7'd325 && y == 170) ||
		(x == 367 && y == 7'd130) || (x == 7'd139 && y == 7'd244) || (x == 7'd624 && y == 315) ||
		(x == 7'd21 && y == 357) || (x == 7'd538 && y == 7'd379) || (x == 585 && y == 301) ||
		(x == 7'd544 && y == 7'd211) || (x == 374 && y == 484) || (x == 342 && y == 379) ||
		(x == 7'd637 && y == 7'd504) || (x == 498 && y == 7'd397) || (x == 198 && y == 640) ||
		(x == 7'd4 && y == 7'd638) || (x == 71 && y == 7'd51) || (x == 7'd252 && y == 7'd575) ||
		(x == 7'd379 && y == 7'd594) || (x == 7'd207 && y == 89) || (x == 7'd57 && y == 7'd16) ||
		(x == 478 && y == 181) || (x == 272 && y == 461) || (x == 7'd374 && y == 7'd446) ||
		(x == 7'd331 && y == 171) || (x == 412 && y == 524) || (x == 7'd532 && y == 7'd523) ||
		(x == 7'd240 && y == 7'd165) || (x == 7'd237 && y == 353) || (x == 7'd25 && y == 636) ||
		(x == 571 && y == 7'd581) || (x == 7'd376 && y == 7'd443) || (x == 7'd572 && y == 7'd89) ||
		(x == 351 && y == 493) || (x == 7'd517 && y == 7'd509) || (x == 7'd232 && y == 7'd497) ||
		(x == 421 && y == 436) || (x == 7'd585 && y == 7'd77) || (x == 506 && y == 382) ||
		(x == 7'd426 && y == 7'd267) || (x == 7'd4 && y == 7'd585) || (x == 636 && y == 608) ||
		(x == 7'd402 && y == 7'd559) || (x == 7'd12 && y == 7'd427) || (x == 7'd578 && y == 273) ||
		(x == 7'd594 && y == 7'd625) || (x == 220 && y == 392) || (x == 90 && y == 7'd497) ||
		(x == 570 && y == 302) || (x == 174 && y == 7'd340) || (x == 385 && y == 7'd149) ||
		(x == 7'd448 && y == 300) || (x == 7'd300 && y == 544) || (x == 377 && y == 7'd509) ||
		(x == 7'd351 && y == 7'd236) || (x == 7'd208 && y == 527) || (x == 593 && y == 286) ||
		(x == 83 && y == 7'd346) || (x == 7'd467 && y == 7'd358) || (x == 7'd535 && y == 272) ||
		(x == 7'd388 && y == 28) || (x == 396 && y == 7'd290) || (x == 476 && y == 7'd132) ||
		(x == 572 && y == 7'd326) || (x == 472 && y == 308) || (x == 7'd428 && y == 83) ||
		(x == 7'd492 && y == 7'd145) || (x == 7'd331 && y == 308) || (x == 7'd295 && y == 7'd470) ||
		(x == 291 && y == 7'd321) || (x == 81 && y == 7'd242) || (x == 7'd216 && y == 7'd41) ||
		(x == 609 && y == 369) || (x == 365 && y == 7'd321) || (x == 611 && y == 7'd405) ||
		(x == 419 && y == 7'd434) || (x == 615 && y == 7'd517) || (x == 16 && y == 7'd0) ||
		(x == 7'd509 && y == 200) || (x == 7'd114 && y == 399) || (x == 616 && y == 7'd590) ||
		(x == 7'd571 && y == 7'd376) || (x == 619 && y == 510) || (x == 533 && y == 460) ||
		(x == 86 && y == 7'd105) || (x == 430 && y == 7'd173) || (x == 7'd462 && y == 7'd345) ||
		(x == 55 && y == 7'd497) || (x == 7'd194 && y == 7'd435) || (x == 594 && y == 7'd28) ||
		(x == 7'd244 && y == 7'd492) || (x == 7'd631 && y == 7'd544) || (x == 590 && y == 7'd92) ||
		(x == 7'd112 && y == 407) || (x == 7'd259 && y == 7'd174) || (x == 7'd285 && y == 460) ||
		(x == 7'd390 && y == 7'd557) || (x == 7'd415 && y == 153) || (x == 574 && y == 141) ||
		(x == 540 && y == 552) || (x == 7'd31 && y == 7'd379) || (x == 7'd155 && y == 7'd262) ||
		(x == 210 && y == 7'd153) || (x == 7'd62 && y == 171) || (x == 274 && y == 7'd488) ||
		(x == 7'd329 && y == 557) || (x == 7'd217 && y == 7'd527) || (x == 7'd380 && y == 7'd615) ||
		(x == 7'd325 && y == 7'd228) || (x == 638 && y == 458) || (x == 361 && y == 7'd73) ||
		(x == 454 && y == 7'd269) || (x == 559 && y == 7'd206) || (x == 276 && y == 600) ||
		(x == 7'd596 && y == 7'd555) || (x == 203 && y == 178) || (x == 7'd200 && y == 474) ||
		(x == 7'd605 && y == 7'd137) || (x == 336 && y == 7'd609) || (x == 7'd528 && y == 7'd319) ||
		(x == 185 && y == 502) || (x == 7'd476 && y == 313) || (x == 7'd193 && y == 39) ||
		(x == 7'd28 && y == 7'd336) || (x == 7'd311 && y == 7'd384) || (x == 7'd382 && y == 7'd537) ||
		(x == 7'd603 && y == 7'd636) || (x == 268 && y == 7'd524) || (x == 7'd62 && y == 7'd374) ||
		(x == 231 && y == 7'd478) || (x == 7'd3 && y == 126) || (x == 7'd238 && y == 324) ||
		(x == 7'd582 && y == 7'd133) || (x == 385 && y == 7'd72) || (x == 40 && y == 7'd503) ||
		(x == 7'd127 && y == 7'd582) || (x == 7'd275 && y == 7'd494) || (x == 594 && y == 7'd35) ||
		(x == 7'd355 && y == 195) || (x == 551 && y == 7'd147) || (x == 601 && y == 594) ||
		(x == 606 && y == 498) || (x == 7'd498 && y == 7'd473) || (x == 7'd154 && y == 453) ||
		(x == 7'd304 && y == 7'd363) || (x == 7'd627 && y == 7'd142) || (x == 7'd579 && y == 7'd187) ||
		(x == 81 && y == 7'd286) || (x == 502 && y == 545) || (x == 7'd639 && y == 230) ||
		(x == 7'd173 && y == 408) || (x == 7'd474 && y == 117) || (x == 7'd574 && y == 7'd448) ||
		(x == 7'd260 && y == 7'd438) || (x == 7'd187 && y == 516) || (x == 7'd351 && y == 7'd362) ||
		(x == 376 && y == 588) || (x == 7'd443 && y == 7'd288) || (x == 634 && y == 7'd25) ||
		(x == 7'd113 && y == 7'd544) || (x == 186 && y == 7'd39) || (x == 7'd534 && y == 68) ||
		(x == 7'd610 && y == 476) || (x == 7'd200 && y == 7'd296) || (x == 287 && y == 7'd399) ||
		(x == 7'd543 && y == 7'd171) || (x == 503 && y == 275) || (x == 7'd236 && y == 361) ||
		(x == 417 && y == 7'd373) || (x == 7'd590 && y == 465) || (x == 7'd123 && y == 7'd442) ||
		(x == 599 && y == 240) || (x == 7'd631 && y == 606) || (x == 7'd302 && y == 217) ||
		(x == 628 && y == 7'd485) || (x == 7'd355 && y == 637) || (x == 3 && y == 7'd183) ||
		(x == 7'd77 && y == 7'd592) || (x == 7'd64 && y == 365) || (x == 7'd202 && y == 7'd42) ||
		(x == 7'd624 && y == 7'd520) || (x == 7'd520 && y == 7'd80) || (x == 7'd544 && y == 7'd141) ||
		(x == 223 && y == 7'd560) || (x == 392 && y == 293) || (x == 7'd243 && y == 7'd312) ||
		(x == 613 && y == 166) || (x == 7'd180 && y == 477) || (x == 7'd553 && y == 7'd376) ||
		(x == 7'd216 && y == 306) || (x == 83 && y == 7'd68) || (x == 7'd574 && y == 7'd87) ||
		(x == 7'd500 && y == 7'd547) || (x == 112 && y == 7'd259) || (x == 7'd129 && y == 510) ||
		(x == 279 && y == 517) || (x == 435 && y == 294) || (x == 41 && y == 7'd178) ||
		(x == 171 && y == 136) || (x == 7'd151 && y == 7'd462) || (x == 517 && y == 7'd1) ||
		(x == 283 && y == 7'd194) || (x == 7'd547 && y == 407) || (x == 396 && y == 7'd458) ||
		(x == 7'd67 && y == 176) || (x == 106 && y == 7'd277) || (x == 325 && y == 7'd635) ||
		(x == 408 && y == 619) || (x == 586 && y == 544) || (x == 422 && y == 357) ||
		(x == 7'd251 && y == 7'd133) || (x == 7'd519 && y == 7'd272) || (x == 589 && y == 7'd528) ||
		(x == 240 && y == 7'd44) || (x == 7'd371 && y == 7'd479) || (x == 132 && y == 506) ||
		(x == 7'd320 && y == 7'd498) || (x == 7'd358 && y == 7'd459) || (x == 452 && y == 7'd134) ||
		(x == 7'd251 && y == 7'd401) || (x == 7'd451 && y == 80) || (x == 595 && y == 389) ||
		(x == 7'd615 && y == 7'd256) || (x == 600 && y == 186) || (x == 526 && y == 433) ||
		(x == 7'd407 && y == 529) || (x == 7'd19 && y == 632) || (x == 7'd432 && y == 7'd388) ||
		(x == 630 && y == 407) || (x == 157 && y == 488) || (x == 7'd541 && y == 210) ||
		(x == 255 && y == 153) || (x == 328 && y == 356) || (x == 7'd394 && y == 7'd241) ||
		(x == 7'd129 && y == 177) || (x == 508 && y == 633) || (x == 7'd123 && y == 7'd227) ||
		(x == 7'd517 && y == 7'd461) || (x == 519 && y == 582) || (x == 133 && y == 7'd616) ||
		(x == 257 && y == 315) || (x == 383 && y == 379) || (x == 16 && y == 7'd295) ||
		(x == 312 && y == 460) || (x == 7'd5 && y == 7'd634) || (x == 204 && y == 7'd135) ||
		(x == 7'd146 && y == 7'd198) || (x == 7'd563 && y == 7'd190) || (x == 127 && y == 7'd619) ||
		(x == 7'd113 && y == 129) || (x == 7'd577 && y == 137) || (x == 48 && y == 7'd528) ||
		(x == 49 && y == 7'd518) || (x == 7'd167 && y == 7'd112) || (x == 7'd159 && y == 7'd363) ||
		(x == 254 && y == 172) || (x == 615 && y == 7'd204) || (x == 7'd392 && y == 592) ||
		(x == 7'd230 && y == 519) || (x == 7'd487 && y == 7'd158) || (x == 243 && y == 373) ||
		(x == 138 && y == 503) || (x == 341 && y == 374) || (x == 381 && y == 7'd34) ||
		(x == 141 && y == 7'd554) || (x == 7'd243 && y == 573) || (x == 7'd580 && y == 7'd37) ||
		(x == 309 && y == 607) || (x == 7'd227 && y == 7'd274) || (x == 7'd347 && y == 7'd165) ||
		(x == 7'd537 && y == 7'd180) || (x == 7'd420 && y == 7'd214) || (x == 7'd25 && y == 388) ||
		(x == 7'd629 && y == 7'd606) || (x == 7'd359 && y == 7'd497) || (x == 7'd597 && y == 7'd174) ||
		(x == 195 && y == 7'd192) || (x == 283 && y == 256) || (x == 7'd164 && y == 7'd500) ||
		(x == 7'd87 && y == 184) || (x == 170 && y == 7'd231) || (x == 7'd108 && y == 534) ||
		(x == 7'd293 && y == 7'd531) || (x == 305 && y == 331) || (x == 7'd353 && y == 7'd211) ||
		(x == 285 && y == 593) || (x == 317 && y == 7'd162) || (x == 485 && y == 235) ||
		(x == 530 && y == 7'd67) || (x == 381 && y == 7'd59) || (x == 7'd202 && y == 7'd173) ||
		(x == 554 && y == 600) || (x == 7'd406 && y == 7'd337) || (x == 201 && y == 7'd45) ||
		(x == 7'd298 && y == 7'd393) || (x == 94 && y == 7'd162) || (x == 348 && y == 7'd576) ||
		(x == 7'd567 && y == 7'd457) || (x == 7'd559 && y == 305) || (x == 7'd452 && y == 7'd254) ||
		(x == 7'd633 && y == 7'd59) || (x == 7'd253 && y == 54) || (x == 544 && y == 7'd542) ||
		(x == 7'd329 && y == 521) || (x == 477 && y == 576) || (x == 518 && y == 7'd183) ||
		(x == 7'd152 && y == 617) || (x == 7'd351 && y == 510) || (x == 7'd391 && y == 7'd556) ||
		(x == 625 && y == 202) || (x == 195 && y == 7'd52) || (x == 7'd468 && y == 4) ||
		(x == 51 && y == 7'd131) || (x == 632 && y == 369) || (x == 593 && y == 7'd566) ||
		(x == 7'd300 && y == 499) || (x == 7'd453 && y == 7'd370) || (x == 7'd216 && y == 419) ||
		(x == 476 && y == 163) || (x == 7'd626 && y == 7'd139) || (x == 7'd8 && y == 7'd621) ||
		(x == 7'd9 && y == 571) || (x == 334 && y == 7'd372) || (x == 7'd351 && y == 7'd11) ||
		(x == 7'd15 && y == 7'd366) || (x == 94 && y == 7'd521) || (x == 7'd545 && y == 7'd363) ||
		(x == 442 && y == 449) || (x == 457 && y == 7'd595) || (x == 7'd245 && y == 7'd546) ||
		(x == 7'd535 && y == 188) || (x == 48 && y == 7'd155) || (x == 7'd203 && y == 7'd306) ||
		(x == 257 && y == 7'd185) || (x == 7'd250 && y == 551) || (x == 7'd573 && y == 245) ||
		(x == 7'd438 && y == 547) || (x == 7'd246 && y == 61) || (x == 7'd465 && y == 7'd538) ||
		(x == 7'd17 && y == 55) || (x == 7'd133 && y == 7'd536) || (x == 447 && y == 167) ||
		(x == 7'd593 && y == 209) || (x == 506 && y == 7'd473) || (x == 255 && y == 7'd393) ||
		(x == 7'd576 && y == 7'd83) || (x == 424 && y == 629) || (x == 624 && y == 7'd577) ||
		(x == 7'd411 && y == 315) || (x == 7'd242 && y == 315) || (x == 550 && y == 259) ||
		(x == 7'd522 && y == 7'd599) || (x == 7'd386 && y == 7'd5) || (x == 203 && y == 241) ||
		(x == 7'd12 && y == 7'd571) || (x == 7'd512 && y == 413) || (x == 171 && y == 7'd6) ||
		(x == 7'd192 && y == 562) || (x == 7'd588 && y == 409) || (x == 7'd323 && y == 7'd560) ||
		(x == 185 && y == 7'd436) || (x == 7'd227 && y == 7'd554) || (x == 7'd99 && y == 302) ||
		(x == 442 && y == 595) || (x == 7'd403 && y == 527) || (x == 323 && y == 639) ||
		(x == 7'd595 && y == 7'd512) || (x == 7'd410 && y == 7'd414) || (x == 16 && y == 7'd527) ||
		(x == 425 && y == 222) || (x == 240 && y == 484) || (x == 7'd502 && y == 609) ||
		(x == 295 && y == 266) || (x == 425 && y == 327) || (x == 7'd577 && y == 7'd541) ||
		(x == 7'd633 && y == 7'd296) || (x == 540 && y == 288) || (x == 167 && y == 193) ||
		(x == 217 && y == 514) || (x == 7'd90 && y == 590) || (x == 334 && y == 7'd344) ||
		(x == 426 && y == 372) || (x == 359 && y == 334) || (x == 149 && y == 7'd445) ||
		(x == 350 && y == 7'd301) || (x == 7'd71 && y == 322) || (x == 7'd566 && y == 130) ||
		(x == 39 && y == 7'd243) || (x == 7'd597 && y == 7'd131) || (x == 7'd35 && y == 97) ||
		(x == 7'd189 && y == 171) || (x == 7'd17 && y == 7'd56) || (x == 7'd285 && y == 589) ||
		(x == 240 && y == 575) || (x == 7'd615 && y == 161) || (x == 633 && y == 504) ||
		(x == 7'd159 && y == 625) || (x == 580 && y == 383) || (x == 7'd342 && y == 7'd259) ||
		(x == 206 && y == 7'd74) || (x == 600 && y == 7'd485) || (x == 7'd146 && y == 7'd160) ||
		(x == 7'd233 && y == 7'd102) || (x == 7'd606 && y == 374) || (x == 7'd183 && y == 7'd276) ||
		(x == 7'd232 && y == 7'd610) || (x == 7'd522 && y == 7'd301) || (x == 162 && y == 436) ||
		(x == 272 && y == 381) || (x == 250 && y == 625) || (x == 7'd220 && y == 7'd525) ||
		(x == 7'd298 && y == 7'd102) || (x == 7'd294 && y == 15) || (x == 180 && y == 7'd203) ||
		(x == 132 && y == 7'd226) || (x == 205 && y == 288) || (x == 7'd358 && y == 7'd506) ||
		(x == 7'd272 && y == 34) || (x == 7'd286 && y == 7'd0) || (x == 632 && y == 305) ||
		(x == 181 && y == 308) || (x == 310 && y == 7'd556) || (x == 7'd393 && y == 7'd377) ||
		(x == 7'd188 && y == 7'd230) || (x == 7'd407 && y == 7'd306) || (x == 189 && y == 7'd189) ||
		(x == 7'd311 && y == 7'd614) || (x == 381 && y == 570) || (x == 7'd478 && y == 7'd493) ||
		(x == 7'd432 && y == 7'd164) || (x == 559 && y == 632) || (x == 7'd508 && y == 483) ||
		(x == 7'd273 && y == 7'd621) || (x == 396 && y == 351) || (x == 7'd144 && y == 7'd281) ||
		(x == 273 && y == 7'd41) || (x == 501 && y == 331) || (x == 127 && y == 44) ||
		(x == 447 && y == 7'd422) || (x == 70 && y == 122) || (x == 7'd638 && y == 7'd75) ||
		(x == 310 && y == 7'd375) || (x == 208 && y == 7'd30) || (x == 7'd415 && y == 1) ||
		(x == 394 && y == 7'd443) || (x == 7'd586 && y == 169) || (x == 628 && y == 7'd491) ||
		(x == 219 && y == 163) || (x == 7'd210 && y == 152) || (x == 591 && y == 499) ||
		(x == 7'd455 && y == 7'd459) || (x == 213 && y == 7'd453) || (x == 134 && y == 7'd363) ||
		(x == 76 && y == 7'd473) || (x == 380 && y == 283) || (x == 113 && y == 7'd420) ||
		(x == 7'd192 && y == 7'd261) || (x == 7'd222 && y == 7'd396) || (x == 288 && y == 7'd399) ||
		(x == 7'd337 && y == 452) || (x == 7'd305 && y == 7'd145) || (x == 7'd496 && y == 95) ||
		(x == 7'd535 && y == 7'd522) || (x == 7'd58 && y == 440) || (x == 7'd82 && y == 7'd331) ||
		(x == 146 && y == 208) || (x == 7'd377 && y == 7'd100) || (x == 7'd131 && y == 466) ||
		(x == 432 && y == 621) || (x == 7'd349 && y == 7'd437) || (x == 7'd409 && y == 7'd557) ||
		(x == 461 && y == 189) || (x == 437 && y == 222) || (x == 630 && y == 7'd507) ||
		(x == 528 && y == 7'd77) || (x == 7'd141 && y == 7'd40) || (x == 338 && y == 7'd73) ||
		(x == 390 && y == 323) || (x == 7'd635 && y == 7'd118) || (x == 7'd51 && y == 298) ||
		(x == 7'd449 && y == 7'd138) || (x == 7'd259 && y == 7'd330) || (x == 7'd312 && y == 67) ||
		(x == 67 && y == 7'd70) || (x == 630 && y == 7'd319) || (x == 7'd76 && y == 7'd285) ||
		(x == 115 && y == 7'd189) || (x == 7'd417 && y == 7'd192) || (x == 406 && y == 617) ||
		(x == 7'd148 && y == 7'd285) || (x == 447 && y == 7'd390) || (x == 7'd319 && y == 7'd371) ||
		(x == 7'd140 && y == 7'd318) || (x == 593 && y == 7'd245) || (x == 614 && y == 7'd605) ||
		(x == 243 && y == 525) || (x == 7'd220 && y == 7'd430) || (x == 7'd126 && y == 272) ||
		(x == 7'd606 && y == 303) || (x == 7'd313 && y == 581) || (x == 7'd173 && y == 330) ||
		(x == 7'd200 && y == 7'd42) || (x == 7'd571 && y == 7'd388) || (x == 7 && y == 7'd577) ||
		(x == 530 && y == 474) || (x == 514 && y == 636) || (x == 138 && y == 7'd502) ||
		(x == 77 && y == 7'd604) || (x == 7'd402 && y == 7'd394) || (x == 7'd397 && y == 7'd150) ||
		(x == 7'd353 && y == 7'd5) || (x == 7'd612 && y == 7'd389) || (x == 148 && y == 7'd163) ||
		(x == 7'd162 && y == 308) || (x == 7'd497 && y == 7'd378) || (x == 7'd316 && y == 381) ||
		(x == 7'd502 && y == 7'd160) || (x == 7'd611 && y == 500) || (x == 381 && y == 7'd241) ||
		(x == 623 && y == 267) || (x == 7'd327 && y == 7'd16) || (x == 157 && y == 614) ||
		(x == 7'd560 && y == 7'd258) || (x == 7'd463 && y == 7'd253) || (x == 530 && y == 129) ||
		(x == 176 && y == 129) || (x == 150 && y == 258) || (x == 7'd310 && y == 7'd144) ||
		(x == 7'd10 && y == 138) || (x == 7'd452 && y == 7'd156) || (x == 7'd221 && y == 7'd397) ||
		(x == 480 && y == 7'd322) || (x == 7'd462 && y == 182) || (x == 7'd362 && y == 7'd562) ||
		(x == 7'd538 && y == 243) || (x == 7'd373 && y == 86) || (x == 7'd479 && y == 527) ||
		(x == 7'd573 && y == 509) || (x == 7'd499 && y == 7'd548) || (x == 555 && y == 7'd464) ||
		(x == 496 && y == 174) || (x == 7'd515 && y == 151) || (x == 7'd357 && y == 7'd241) ||
		(x == 284 && y == 7'd544) || (x == 326 && y == 7'd416) || (x == 261 && y == 600) ||
		(x == 7'd63 && y == 603) || (x == 7'd74 && y == 370) || (x == 593 && y == 571) ||
		(x == 7'd345 && y == 494) || (x == 604 && y == 633) || (x == 7'd466 && y == 7'd569) ||
		(x == 7'd277 && y == 7'd437) || (x == 7'd251 && y == 7'd229) || (x == 7'd114 && y == 7'd288) ||
		(x == 132 && y == 583) || (x == 321 && y == 401) || (x == 576 && y == 7'd13) ||
		(x == 630 && y == 544) || (x == 7'd445 && y == 205) || (x == 395 && y == 640) ||
		(x == 354 && y == 620) || (x == 273 && y == 7'd576) || (x == 433 && y == 343) ||
		(x == 7'd186 && y == 406) || (x == 7'd319 && y == 7'd423) || (x == 7'd227 && y == 7'd638) ||
		(x == 7'd154 && y == 7'd135) || (x == 457 && y == 7'd525) || (x == 211 && y == 7'd406) ||
		(x == 164 && y == 316) || (x == 7'd617 && y == 133) || (x == 7'd475 && y == 446) ||
		(x == 7'd349 && y == 289) || (x == 281 && y == 232) || (x == 213 && y == 315) ||
		(x == 7'd189 && y == 538) || (x == 448 && y == 602) || (x == 7'd248 && y == 7'd229) ||
		(x == 235 && y == 502) || (x == 337 && y == 7'd537) || (x == 185 && y == 448) ||
		(x == 435 && y == 340) || (x == 7'd107 && y == 179) || (x == 7'd146 && y == 7'd211) ||
		(x == 7'd463 && y == 405) || (x == 7'd236 && y == 635) || (x == 35 && y == 7'd131) ||
		(x == 7'd405 && y == 7'd518) || (x == 631 && y == 7'd512) || (x == 7'd65 && y == 7'd133) ||
		(x == 7'd391 && y == 7'd395) || (x == 420 && y == 502) || (x == 637 && y == 446) ||
		(x == 450 && y == 7'd189) || (x == 7'd619 && y == 7'd228) || (x == 482 && y == 388) ||
		(x == 7'd346 && y == 593) || (x == 406 && y == 7'd1) || (x == 398 && y == 7'd508) ||
		(x == 7'd328 && y == 41) || (x == 7'd431 && y == 309) || (x == 72 && y == 7'd617) ||
		(x == 129 && y == 628) || (x == 312 && y == 363) || (x == 7'd288 && y == 7'd502) ||
		(x == 533 && y == 343) || (x == 7'd393 && y == 21) || (x == 7'd478 && y == 614) ||
		(x == 7'd423 && y == 547) || (x == 7'd300 && y == 376) || (x == 207 && y == 552) ||
		(x == 7'd21 && y == 339) || (x == 4 && y == 66) || (x == 7'd228 && y == 7'd171) ||
		(x == 187 && y == 7'd59) || (x == 7'd272 && y == 7'd524) || (x == 293 && y == 288) ||
		(x == 7'd236 && y == 7'd561) || (x == 434 && y == 7'd606) || (x == 582 && y == 7'd92) ||
		(x == 7'd453 && y == 605) || (x == 193 && y == 352) || (x == 7'd93 && y == 289) ||
		(x == 537 && y == 383) || (x == 7'd247 && y == 527) || (x == 263 && y == 7'd492) ||
		(x == 7'd210 && y == 292) || (x == 7'd316 && y == 308) || (x == 532 && y == 387) ||
		(x == 380 && y == 497) || (x == 7'd23 && y == 7'd262) || (x == 7'd497 && y == 363) ||
		(x == 401 && y == 7'd50) || (x == 184 && y == 7'd289) || (x == 7'd285 && y == 7'd395) ||
		(x == 504 && y == 7'd295) || (x == 163 && y == 7'd30) || (x == 463 && y == 7'd390) ||
		(x == 7'd615 && y == 45) || (x == 253 && y == 7'd478) || (x == 7'd320 && y == 7'd519) ||
		(x == 435 && y == 7'd100) || (x == 7'd66 && y == 7'd561) || (x == 7'd355 && y == 7'd494) ||
		(x == 202 && y == 7'd546) || (x == 7'd576 && y == 7'd398) || (x == 7'd446 && y == 7'd520) ||
		(x == 7'd253 && y == 7'd210) || (x == 350 && y == 472) || (x == 7'd517 && y == 7'd520) ||
		(x == 7'd600 && y == 440) || (x == 515 && y == 559) || (x == 7'd639 && y == 323) ||
		(x == 555 && y == 291) || (x == 7'd321 && y == 7'd96) || (x == 577 && y == 214) ||
		(x == 7'd564 && y == 247) || (x == 7'd558 && y == 548) || (x == 206 && y == 7'd410) ||
		(x == 7'd54 && y == 218) || (x == 342 && y == 7'd571) || (x == 7'd592 && y == 550) ||
		(x == 7'd104 && y == 7'd122) || (x == 7'd446 && y == 7'd131) || (x == 7'd492 && y == 7'd405) ||
		(x == 7'd267 && y == 7'd375) || (x == 7'd483 && y == 7'd636) || (x == 188 && y == 312) ||
		(x == 7'd166 && y == 7'd471) || (x == 7'd519 && y == 42) || (x == 458 && y == 492) ||
		(x == 7'd608 && y == 7'd235) || (x == 7'd578 && y == 7'd422) || (x == 201 && y == 7'd459) ||
		(x == 428 && y == 546) || (x == 7'd458 && y == 7'd132) || (x == 5 && y == 7'd289) ||
		(x == 7'd639 && y == 7'd617) || (x == 385 && y == 7'd533) || (x == 7'd447 && y == 7'd133) ||
		(x == 535 && y == 7'd33) || (x == 522 && y == 636) || (x == 7'd458 && y == 7'd491) ||
		(x == 7'd484 && y == 326) || (x == 7'd111 && y == 7'd389) || (x == 7'd581 && y == 7'd391) ||
		(x == 7'd598 && y == 7'd478) || (x == 563 && y == 7'd461) || (x == 7'd379 && y == 7'd339) ||
		(x == 7'd458 && y == 7'd529) || (x == 7'd335 && y == 7'd113) || (x == 337 && y == 530) ||
		(x == 246 && y == 7'd505) || (x == 522 && y == 203) || (x == 401 && y == 587) ||
		(x == 7'd403 && y == 7'd207) || (x == 524 && y == 267) || (x == 192 && y == 7'd560) ||
		(x == 281 && y == 552) || (x == 7'd237 && y == 588) || (x == 7'd6 && y == 7'd163) ||
		(x == 276 && y == 466) || (x == 559 && y == 334) || (x == 7'd237 && y == 7'd428) ||
		(x == 473 && y == 566) || (x == 7'd261 && y == 7'd332) || (x == 7'd258 && y == 7'd71) ||
		(x == 403 && y == 7'd504) || (x == 7'd108 && y == 7'd560) || (x == 58 && y == 7'd352) ||
		(x == 7'd337 && y == 393) || (x == 535 && y == 7'd560) || (x == 556 && y == 7'd622) ||
		(x == 102 && y == 76) || (x == 611 && y == 7'd148) || (x == 7'd298 && y == 7'd398) ||
		(x == 7'd500 && y == 7'd164) || (x == 577 && y == 593) || (x == 134 && y == 581) ||
		(x == 542 && y == 7'd415) || (x == 7'd541 && y == 54) || (x == 7'd625 && y == 7'd581) ||
		(x == 7'd132 && y == 7'd619) || (x == 7'd90 && y == 241) || (x == 7'd286 && y == 483) ||
		(x == 623 && y == 7'd80) || (x == 7'd180 && y == 7'd310) || (x == 7'd183 && y == 7'd584) ||
		(x == 7'd514 && y == 7'd361) || (x == 7'd355 && y == 200) || (x == 176 && y == 560) ||
		(x == 7'd568 && y == 633) || (x == 627 && y == 431) || (x == 565 && y == 7'd10) ||
		(x == 7'd296 && y == 7'd261) || (x == 7'd320 && y == 7'd373) || (x == 7'd455 && y == 125) ||
		(x == 238 && y == 7'd611) || (x == 7'd353 && y == 7'd286) || (x == 412 && y == 7'd19) ||
		(x == 7'd195 && y == 7'd206) || (x == 7'd215 && y == 358) || (x == 422 && y == 7'd445) ||
		(x == 7'd55 && y == 169) || (x == 7'd145 && y == 7'd41) || (x == 7'd198 && y == 188) ||
		(x == 7'd318 && y == 526) || (x == 7'd637 && y == 7'd247) || (x == 7'd329 && y == 7'd235) ||
		(x == 546 && y == 203) || (x == 7'd582 && y == 7'd111) || (x == 466 && y == 603) ||
		(x == 74 && y == 7'd309) || (x == 240 && y == 7'd235) || (x == 632 && y == 132) ||
		(x == 7'd321 && y == 7'd216) || (x == 461 && y == 7'd375) || (x == 561 && y == 7'd389) ||
		(x == 7'd315 && y == 7'd500) || (x == 173 && y == 7'd84) || (x == 7'd557 && y == 497) ||
		(x == 310 && y == 7'd549) || (x == 7'd523 && y == 7'd216) || (x == 7'd429 && y == 285) ||
		(x == 7'd448 && y == 224) || (x == 469 && y == 7'd40) || (x == 7'd374 && y == 7'd542) ||
		(x == 517 && y == 134) || (x == 241 && y == 325) || (x == 7'd223 && y == 404) ||
		(x == 7'd320 && y == 426) || (x == 7'd281 && y == 243) || (x == 7'd472 && y == 307) ||
		(x == 7'd481 && y == 7'd364) || (x == 7'd358 && y == 7'd626) || (x == 130 && y == 161) ||
		(x == 380 && y == 622) || (x == 291 && y == 7'd33) || (x == 357 && y == 299) ||
		(x == 7'd362 && y == 7'd480) || (x == 7'd234 && y == 116) || (x == 7'd274 && y == 348) ||
		(x == 524 && y == 7'd172) || (x == 7'd407 && y == 7'd204) || (x == 7'd320 && y == 189) ||
		(x == 544 && y == 531) || (x == 7'd72 && y == 318) || (x == 7'd536 && y == 7'd558) ||
		(x == 546 && y == 7'd610) || (x == 7'd301 && y == 7'd139) || (x == 7'd354 && y == 7'd400) ||
		(x == 7'd624 && y == 7'd182) || (x == 455 && y == 7'd454) || (x == 7'd250 && y == 7'd356) ||
		(x == 506 && y == 7'd113) || (x == 7'd418 && y == 7'd275) || (x == 566 && y == 413) ||
		(x == 7'd230 && y == 7'd428) || (x == 7'd461 && y == 7'd403) || (x == 7'd207 && y == 7'd626) ||
		(x == 537 && y == 7'd155) || (x == 320 && y == 269) || (x == 547 && y == 7'd456) ||
		(x == 118 && y == 7'd262) || (x == 461 && y == 538) || (x == 7'd552 && y == 214) ||
		(x == 366 && y == 7'd125) || (x == 7'd149 && y == 7'd455) || (x == 7'd217 && y == 438) ||
		(x == 424 && y == 7'd194) || (x == 7'd443 && y == 7'd274) || (x == 7'd228 && y == 7'd131) ||
		(x == 7'd346 && y == 476) || (x == 7'd312 && y == 7'd148) || (x == 7'd519 && y == 7'd419) ||
		(x == 321 && y == 259) || (x == 7'd121 && y == 5) || (x == 508 && y == 7'd129) ||
		(x == 561 && y == 7'd451) || (x == 7'd193 && y == 7'd498) || (x == 7'd498 && y == 7'd308) ||
		(x == 15 && y == 7'd469) || (x == 202 && y == 386) || (x == 7'd464 && y == 7'd239) ||
		(x == 7'd393 && y == 257) || (x == 235 && y == 144) || (x == 7'd348 && y == 437) ||
		(x == 7'd344 && y == 7'd164) || (x == 7'd394 && y == 7'd40) || (x == 7'd278 && y == 7'd565) ||
		(x == 7'd518 && y == 7'd143) || (x == 7'd369 && y == 7'd545) || (x == 7'd218 && y == 7'd633) ||
		(x == 7'd497 && y == 7'd348) || (x == 7'd86 && y == 603) || (x == 562 && y == 326) ||
		(x == 614 && y == 7'd399) || (x == 7'd603 && y == 633) || (x == 7'd66 && y == 7'd548) ||
		(x == 7'd479 && y == 639) || (x == 7'd628 && y == 408) || (x == 7'd476 && y == 7'd462) ||
		(x == 7'd80 && y == 521) || (x == 7'd570 && y == 7'd353) || (x == 7'd638 && y == 98) ||
		(x == 418 && y == 7'd471) || (x == 7'd578 && y == 37) || (x == 457 && y == 7'd167) ||
		(x == 11 && y == 7'd425) || (x == 7'd485 && y == 7'd334) || (x == 7'd243 && y == 279) ||
		(x == 7'd162 && y == 7'd38) || (x == 7'd202 && y == 7'd398) || (x == 7'd214 && y == 7'd177) ||
		(x == 123 && y == 7'd543) || (x == 270 && y == 267) || (x == 7'd132 && y == 374) ||
		(x == 7'd169 && y == 7'd520) || (x == 324 && y == 7'd460) || (x == 261 && y == 7'd403) ||
		(x == 7'd421 && y == 7'd271) || (x == 7'd53 && y == 606) || (x == 416 && y == 7'd338) ||
		(x == 197 && y == 7'd359) || (x == 7'd188 && y == 7'd274) || (x == 211 && y == 520) ||
		(x == 7'd262 && y == 420) || (x == 7'd225 && y == 328) || (x == 501 && y == 366) ||
		(x == 7'd307 && y == 13) || (x == 232 && y == 7'd82) || (x == 238 && y == 7'd103) ||
		(x == 548 && y == 7'd589) || (x == 598 && y == 7'd490) || (x == 157 && y == 7'd615) ||
		(x == 7'd143 && y == 227) || (x == 7'd239 && y == 7'd306) || (x == 7'd105 && y == 420) ||
		(x == 7'd41 && y == 7'd11) || (x == 582 && y == 198) || (x == 7'd386 && y == 7'd154) ||
		(x == 575 && y == 7'd8) || (x == 419 && y == 518) || (x == 7'd9 && y == 20) ||
		(x == 351 && y == 622) || (x == 7'd248 && y == 7'd271) || (x == 177 && y == 7'd16) ||
		(x == 7'd250 && y == 7'd258) || (x == 7'd561 && y == 7'd80) || (x == 7'd333 && y == 7'd428) ||
		(x == 7'd615 && y == 7'd335) || (x == 7'd573 && y == 419) || (x == 7'd75 && y == 203) ||
		(x == 7'd442 && y == 445) || (x == 33 && y == 7'd578) || (x == 7'd46 && y == 553) ||
		(x == 243 && y == 7'd14) || (x == 316 && y == 207) || (x == 7'd200 && y == 7'd495) ||
		(x == 407 && y == 475) || (x == 7'd188 && y == 7'd635) || (x == 531 && y == 7'd368) ||
		(x == 7'd371 && y == 7'd320) || (x == 7'd201 && y == 549) || (x == 7'd529 && y == 7'd273) ||
		(x == 69 && y == 7'd607) || (x == 7'd339 && y == 454) || (x == 7'd571 && y == 7'd369) ||
		(x == 198 && y == 542) || (x == 7'd619 && y == 7'd274) || (x == 7'd388 && y == 7'd351) ||
		(x == 199 && y == 253) || (x == 571 && y == 7'd399) || (x == 7'd359 && y == 7'd230) ||
		(x == 7'd293 && y == 7'd600) || (x == 7'd404 && y == 7'd619) || (x == 7'd73 && y == 7'd423) ||
		(x == 435 && y == 519) || (x == 612 && y == 224) || (x == 157 && y == 286) ||
		(x == 7'd536 && y == 7'd176) || (x == 509 && y == 455) || (x == 326 && y == 7'd562) ||
		(x == 7'd515 && y == 318) || (x == 7'd344 && y == 7'd549) || (x == 7'd619 && y == 7'd404) ||
		(x == 7'd148 && y == 7'd300) || (x == 517 && y == 7'd485) || (x == 7'd82 && y == 568) ||
		(x == 214 && y == 239) || (x == 507 && y == 312) || (x == 133 && y == 7'd162) ||
		(x == 7'd325 && y == 7'd296) || (x == 327 && y == 557) || (x == 7'd637 && y == 7'd588) ||
		(x == 7'd247 && y == 7'd523) || (x == 7'd471 && y == 7'd167) || (x == 7'd164 && y == 7'd596) ||
		(x == 391 && y == 7'd526) || (x == 7'd262 && y == 7'd578) || (x == 7'd12 && y == 7'd316) ||
		(x == 7'd326 && y == 616) || (x == 613 && y == 7'd309) || (x == 7'd516 && y == 7'd260) ||
		(x == 7'd523 && y == 65) || (x == 117 && y == 7'd587) || (x == 561 && y == 540) ||
		(x == 518 && y == 7'd161) || (x == 330 && y == 361) || (x == 7'd278 && y == 575) ||
		(x == 7'd479 && y == 409) || (x == 7'd452 && y == 365) || (x == 7'd381 && y == 186) ||
		(x == 7'd198 && y == 7'd260) || (x == 229 && y == 428) || (x == 520 && y == 640) ||
		(x == 321 && y == 7'd619) || (x == 530 && y == 377) || (x == 7'd131 && y == 7'd264) ||
		(x == 7'd195 && y == 308) || (x == 513 && y == 7'd39) || (x == 333 && y == 7'd555) ||
		(x == 7'd414 && y == 7'd617) || (x == 7'd354 && y == 7'd525) || (x == 7'd130 && y == 7'd565) ||
		(x == 7'd492 && y == 529) || (x == 216 && y == 7'd359) || (x == 344 && y == 139) ||
		(x == 7'd232 && y == 636) || (x == 7'd79 && y == 513) || (x == 7'd575 && y == 263) ||
		(x == 7'd407 && y == 462) || (x == 308 && y == 7'd593) || (x == 383 && y == 171) ||
		(x == 615 && y == 7'd562) || (x == 446 && y == 7'd303) || (x == 7'd434 && y == 536) ||
		(x == 7'd370 && y == 7'd124) || (x == 7'd428 && y == 452) || (x == 7'd336 && y == 189) ||
		(x == 150 && y == 134) || (x == 118 && y == 7'd227) || (x == 7'd424 && y == 7'd598) ||
		(x == 7'd62 && y == 226) || (x == 7'd411 && y == 7'd183) || (x == 7'd510 && y == 584) ||
		(x == 7'd7 && y == 7'd431) || (x == 7'd517 && y == 145) || (x == 321 && y == 590) ||
		(x == 7'd460 && y == 7'd483) || (x == 329 && y == 182) || (x == 7'd491 && y == 7'd154) ||
		(x == 7'd621 && y == 7'd88) || (x == 7'd607 && y == 7'd268) || (x == 7'd138 && y == 7'd165) ||
		(x == 7'd586 && y == 478) || (x == 343 && y == 7'd105) || (x == 7'd195 && y == 7'd139) ||
		(x == 7'd209 && y == 324) || (x == 402 && y == 7'd585) || (x == 10 && y == 7'd193) ||
		(x == 386 && y == 318) || (x == 396 && y == 427) || (x == 7'd89 && y == 386) ||
		(x == 7'd136 && y == 7'd567) || (x == 100 && y == 7'd636) || (x == 7'd90 && y == 40) ||
		(x == 7'd507 && y == 7'd515) || (x == 7'd453 && y == 7'd239) || (x == 7'd561 && y == 7'd267) ||
		(x == 7'd175 && y == 7'd393) || (x == 7'd236 && y == 7'd95) || (x == 388 && y == 7'd130) ||
		(x == 7'd248 && y == 362) || (x == 539 && y == 182) || (x == 7'd358 && y == 541) ||
		(x == 7'd530 && y == 7'd619) || (x == 286 && y == 194) || (x == 7'd565 && y == 7'd274) ||
		(x == 7'd352 && y == 7'd518) || (x == 635 && y == 7'd560) || (x == 475 && y == 330) ||
		(x == 7'd122 && y == 519) || (x == 570 && y == 7'd617) || (x == 7'd339 && y == 7'd570) ||
		(x == 7'd79 && y == 621) || (x == 7'd500 && y == 7'd549) || (x == 318 && y == 7'd164) ||
		(x == 187 && y == 233) || (x == 7'd104 && y == 279) || (x == 7'd605 && y == 7'd367) ||
		(x == 7'd371 && y == 7'd347) || (x == 7'd368 && y == 7'd89) || (x == 7'd124 && y == 298) ||
		(x == 7'd535 && y == 556) || (x == 7'd514 && y == 168) || (x == 7'd13 && y == 415) ||
		(x == 502 && y == 611) || (x == 422 && y == 496) || (x == 7'd512 && y == 235) ||
		(x == 7'd209 && y == 7'd338) || (x == 360 && y == 374) || (x == 7'd252 && y == 435) ||
		(x == 7'd599 && y == 7'd143) || (x == 7'd103 && y == 280) || (x == 7'd376 && y == 7'd442) ||
		(x == 326 && y == 233) || (x == 7'd453 && y == 7'd72) || (x == 7'd600 && y == 7'd377) ||
		(x == 7'd378 && y == 7'd314) || (x == 7'd636 && y == 7'd542) || (x == 237 && y == 7'd634) ||
		(x == 242 && y == 408) || (x == 124 && y == 7'd451) || (x == 7'd240 && y == 430) ||
		(x == 263 && y == 196) || (x == 7'd604 && y == 391) || (x == 7'd403 && y == 7'd47) ||
		(x == 441 && y == 227) || (x == 145 && y == 284) || (x == 374 && y == 7'd118) ||
		(x == 7'd59 && y == 198) || (x == 7'd376 && y == 7'd356) || (x == 7'd177 && y == 7'd260) ||
		(x == 396 && y == 208) || (x == 7'd598 && y == 258) || (x == 7'd178 && y == 7'd223) ||
		(x == 7'd137 && y == 556) || (x == 7'd136 && y == 7'd543) || (x == 616 && y == 7'd602) ||
		(x == 7'd54 && y == 7'd403) || (x == 234 && y == 421) || (x == 7'd473 && y == 7'd180) ||
		(x == 379 && y == 7'd167) || (x == 492 && y == 7'd229) || (x == 342 && y == 7'd89) ||
		(x == 7'd191 && y == 325) || (x == 7'd413 && y == 7'd522) || (x == 264 && y == 589) ||
		(x == 7'd346 && y == 7'd11) || (x == 274 && y == 7'd220) || (x == 7'd78 && y == 241) ||
		(x == 7'd344 && y == 174) || (x == 7'd419 && y == 7'd235) || (x == 131 && y == 304) ||
		(x == 7'd491 && y == 356) || (x == 396 && y == 586) || (x == 168 && y == 291) ||
		(x == 7'd532 && y == 7'd279) || (x == 7'd598 && y == 153) || (x == 451 && y == 134) ||
		(x == 7'd493 && y == 7'd45) || (x == 7'd142 && y == 115) || (x == 7'd378 && y == 7'd297) ||
		(x == 473 && y == 561) || (x == 627 && y == 573) || (x == 7'd154 && y == 7'd514) ||
		(x == 484 && y == 7'd619) || (x == 7'd294 && y == 7'd89) || (x == 7'd25 && y == 262) ||
		(x == 446 && y == 567) || (x == 126 && y == 7'd364) || (x == 462 && y == 7'd317) ||
		(x == 588 && y == 7'd480) || (x == 249 && y == 7'd393) || (x == 270 && y == 7'd464) ||
		(x == 7'd185 && y == 7'd498) || (x == 7'd473 && y == 5) || (x == 7'd613 && y == 7'd429) ||
		(x == 7'd479 && y == 551) || (x == 7'd232 && y == 7'd302) || (x == 116 && y == 7'd90) ||
		(x == 7'd336 && y == 7'd378) || (x == 152 && y == 227) || (x == 7'd399 && y == 7'd502) ||
		(x == 140 && y == 7'd523) || (x == 171 && y == 7'd212) || (x == 7'd388 && y == 7'd454) ||
		(x == 7'd640 && y == 254) || (x == 7'd418 && y == 217) || (x == 112 && y == 7'd196) ||
		(x == 369 && y == 594) || (x == 398 && y == 633) || (x == 7'd318 && y == 7'd415) ||
		(x == 7'd20 && y == 82) || (x == 422 && y == 7'd360) || (x == 7'd471 && y == 7'd631) ||
		(x == 7'd500 && y == 7'd314) || (x == 7'd73 && y == 218) || (x == 217 && y == 7'd128) ||
		(x == 152 && y == 424) || (x == 327 && y == 283) || (x == 7'd601 && y == 238) ||
		(x == 7'd191 && y == 7'd195) || (x == 7'd427 && y == 7'd338) || (x == 246 && y == 422) ||
		(x == 7'd168 && y == 7'd519) || (x == 363 && y == 7'd594) || (x == 7'd157 && y == 7'd418) ||
		(x == 130 && y == 7'd549) || (x == 636 && y == 206) || (x == 7'd252 && y == 7'd517) ||
		(x == 7'd380 && y == 7'd272) || (x == 7'd342 && y == 289) || (x == 7'd497 && y == 7'd424) ||
		(x == 7'd227 && y == 7'd106) || (x == 601 && y == 7'd206) || (x == 506 && y == 7'd480) ||
		(x == 7'd568 && y == 550) || (x == 7'd566 && y == 7'd585) || (x == 7'd283 && y == 7'd388) ||
		(x == 238 && y == 264) || (x == 518 && y == 324) || (x == 637 && y == 628) ||
		(x == 7'd62 && y == 7'd98) || (x == 457 && y == 199) || (x == 507 && y == 372) ||
		(x == 571 && y == 256) || (x == 7'd376 && y == 7'd311) || (x == 7'd560 && y == 425) ||
		(x == 522 && y == 487) || (x == 7'd597 && y == 7'd475) || (x == 7'd427 && y == 572) ||
		(x == 366 && y == 7'd112) || (x == 7'd273 && y == 120) || (x == 7'd405 && y == 534) ||
		(x == 7'd582 && y == 7'd570) || (x == 7'd451 && y == 7'd164) || (x == 541 && y == 258) ||
		(x == 7'd514 && y == 142) || (x == 7'd404 && y == 197) || (x == 20 && y == 7'd306) ||
		(x == 7'd605 && y == 48) || (x == 549 && y == 570) || (x == 7'd188 && y == 169) ||
		(x == 534 && y == 7'd112) || (x == 581 && y == 513) || (x == 418 && y == 7'd40) ||
		(x == 246 && y == 635) || (x == 191 && y == 347) || (x == 566 && y == 541) ||
		(x == 7'd586 && y == 7'd439) || (x == 611 && y == 533) || (x == 7'd292 && y == 413) ||
		(x == 429 && y == 171) || (x == 346 && y == 584) || (x == 516 && y == 7'd267) ||
		(x == 431 && y == 431) || (x == 7'd403 && y == 7'd386) || (x == 7'd377 && y == 7'd590) ||
		(x == 7'd578 && y == 524) || (x == 7'd541 && y == 7'd181) || (x == 386 && y == 240) ||
		(x == 7'd398 && y == 7'd217) || (x == 216 && y == 158) || (x == 386 && y == 582) ||
		(x == 7'd302 && y == 7'd508) || (x == 7'd634 && y == 560) || (x == 7'd239 && y == 313) ||
		(x == 336 && y == 7'd79) || (x == 7'd278 && y == 7'd3) || (x == 333 && y == 7'd188) ||
		(x == 558 && y == 7'd285) || (x == 226 && y == 7'd72) || (x == 539 && y == 7'd569) ||
		(x == 19 && y == 7'd163) || (x == 293 && y == 7'd193) || (x == 502 && y == 7'd71) ||
		(x == 7'd249 && y == 7'd591) || (x == 271 && y == 252) || (x == 7'd266 && y == 0) ||
		(x == 7'd319 && y == 193) || (x == 7'd561 && y == 7'd607) || (x == 7'd296 && y == 216) ||
		(x == 621 && y == 456) || (x == 7'd282 && y == 7'd167) || (x == 7'd90 && y == 250) ||
		(x == 7'd572 && y == 576) || (x == 583 && y == 369) || (x == 7'd29 && y == 7'd556) ||
		(x == 7'd158 && y == 7'd608) || (x == 7'd301 && y == 7'd382) || (x == 7'd163 && y == 369) ||
		(x == 7'd336 && y == 169) || (x == 7'd395 && y == 7'd270) || (x == 252 && y == 223) ||
		(x == 7'd14 && y == 359) || (x == 7'd413 && y == 210) || (x == 7'd542 && y == 7'd379) ||
		(x == 7'd295 && y == 355) || (x == 409 && y == 7'd507) || (x == 7'd101 && y == 7'd366) ||
		(x == 395 && y == 7'd171) || (x == 119 && y == 7'd466) || (x == 7'd630 && y == 7'd607) ||
		(x == 7'd497 && y == 7'd504) || (x == 7'd612 && y == 7'd401) || (x == 7'd80 && y == 134) ||
		(x == 564 && y == 7'd184) || (x == 358 && y == 7'd430) || (x == 7'd516 && y == 7'd195) ||
		(x == 7'd330 && y == 7'd399) || (x == 417 && y == 7'd437) || (x == 7'd624 && y == 7'd451) ||
		(x == 7'd136 && y == 7'd378) || (x == 7'd272 && y == 7'd248) || (x == 7'd270 && y == 7'd147) ||
		(x == 7'd263 && y == 7'd398) || (x == 7'd556 && y == 7'd230) || (x == 7'd261 && y == 515) ||
		(x == 7'd487 && y == 7'd368) || (x == 7'd601 && y == 7'd163) || (x == 7'd324 && y == 7'd304) ||
		(x == 7'd557 && y == 225) || (x == 359 && y == 7'd311) || (x == 7'd572 && y == 414) ||
		(x == 395 && y == 549) || (x == 7'd207 && y == 7'd403) || (x == 129 && y == 7'd387) ||
		(x == 99 && y == 7'd488) || (x == 617 && y == 635) || (x == 165 && y == 419) ||
		(x == 316 && y == 362) || (x == 339 && y == 7'd385) || (x == 196 && y == 345) ||
		(x == 7'd109 && y == 626) || (x == 570 && y == 7'd199) || (x == 19 && y == 32) ||
		(x == 7'd125 && y == 143) || (x == 409 && y == 7'd206) || (x == 472 && y == 237) ||
		(x == 250 && y == 570) || (x == 7'd607 && y == 7'd527) || (x == 189 && y == 7'd344) ||
		(x == 501 && y == 622) || (x == 7'd148 && y == 223) || (x == 212 && y == 308) ||
		(x == 8 && y == 7'd556) || (x == 295 && y == 357) || (x == 7'd229 && y == 7'd331) ||
		(x == 464 && y == 539) || (x == 569 && y == 7'd557) || (x == 7'd135 && y == 7'd250) ||
		(x == 7'd591 && y == 7'd341) || (x == 7'd196 && y == 7'd584) || (x == 7'd329 && y == 55) ||
		(x == 7'd482 && y == 547) || (x == 592 && y == 7'd246) || (x == 560 && y == 435) ||
		(x == 445 && y == 7'd484) || (x == 7'd438 && y == 7'd72) || (x == 592 && y == 7'd230) ||
		(x == 7'd309 && y == 7'd76) || (x == 609 && y == 511) || (x == 309 && y == 7'd92) ||
		(x == 254 && y == 191) || (x == 7'd130 && y == 299) || (x == 7'd63 && y == 328) ||
		(x == 7'd324 && y == 7'd313) || (x == 7'd611 && y == 7'd568) || (x == 333 && y == 628) ||
		(x == 7'd395 && y == 7'd594) || (x == 7'd156 && y == 276) || (x == 7'd469 && y == 7'd212) ||
		(x == 592 && y == 269) || (x == 7'd625 && y == 245) || (x == 7'd334 && y == 7'd539) ||
		(x == 118 && y == 7'd519) || (x == 14 && y == 7'd471) || (x == 32 && y == 119) ||
		(x == 7'd139 && y == 7'd549) || (x == 7'd252 && y == 7'd424) || (x == 7'd235 && y == 7'd553) ||
		(x == 623 && y == 7'd286) || (x == 7'd422 && y == 7'd458) || (x == 284 && y == 7'd177) ||
		(x == 7'd361 && y == 7'd275) || (x == 419 && y == 589) || (x == 7'd116 && y == 399) ||
		(x == 571 && y == 7'd168) || (x == 595 && y == 7'd312) || (x == 7'd530 && y == 7'd398) ||
		(x == 7'd381 && y == 605) || (x == 465 && y == 7'd538) || (x == 223 && y == 612) ||
		(x == 7'd579 && y == 7'd340) || (x == 195 && y == 7'd452) || (x == 7'd158 && y == 7'd523) ||
		(x == 7'd608 && y == 465) || (x == 7'd499 && y == 7'd449) || (x == 7'd115 && y == 7'd523) ||
		(x == 7'd509 && y == 7'd321) || (x == 7'd287 && y == 364) || (x == 265 && y == 7'd598) ||
		(x == 7'd292 && y == 440) || (x == 7'd372 && y == 7'd199) || (x == 291 && y == 7'd19) ||
		(x == 7'd312 && y == 245) || (x == 7'd46 && y == 7'd7) || (x == 184 && y == 7'd213) ||
		(x == 7'd521 && y == 7'd430) || (x == 597 && y == 7'd254) || (x == 325 && y == 380) ||
		(x == 7'd596 && y == 495) || (x == 292 && y == 183) || (x == 7'd448 && y == 7'd341) ||
		(x == 282 && y == 234) || (x == 337 && y == 7'd587) || (x == 588 && y == 519) ||
		(x == 19 && y == 7'd504) || (x == 122 && y == 7'd588) || (x == 162 && y == 7'd313) ||
		(x == 7'd467 && y == 7'd114) || (x == 7'd416 && y == 169) || (x == 124 && y == 7'd411) ||
		(x == 7'd550 && y == 7'd389) || (x == 638 && y == 233) || (x == 7'd622 && y == 7'd275) ||
		(x == 7'd427 && y == 7'd138) || (x == 518 && y == 7'd261) || (x == 7'd474 && y == 7'd144) ||
		(x == 12 && y == 84) || (x == 7'd80 && y == 7'd123) || (x == 7'd501 && y == 7'd349) ||
		(x == 7'd531 && y == 384) || (x == 7'd527 && y == 7'd2) || (x == 7'd13 && y == 7'd473) ||
		(x == 7'd29 && y == 7'd293) || (x == 7'd551 && y == 7'd374) || (x == 7'd105 && y == 7'd175) ||
		(x == 7'd425 && y == 7'd214) || (x == 579 && y == 7'd190) || (x == 7'd638 && y == 18) ||
		(x == 7'd194 && y == 7'd336) || (x == 7'd80 && y == 232) || (x == 7'd565 && y == 7'd296) ||
		(x == 7'd544 && y == 7'd579) || (x == 7'd363 && y == 7'd539) || (x == 7'd134 && y == 7'd397) ||
		(x == 7'd176 && y == 7'd588) || (x == 7'd447 && y == 7'd396) || (x == 7'd619 && y == 7'd502) ||
		(x == 7'd366 && y == 7'd143) || (x == 216 && y == 586) || (x == 7'd338 && y == 7'd455) ||
		(x == 379 && y == 7'd593) || (x == 7'd526 && y == 7'd426) || (x == 7'd589 && y == 7'd90) ||
		(x == 7'd390 && y == 7'd476) || (x == 7'd231 && y == 7'd239) || (x == 7'd284 && y == 7'd256) ||
		(x == 149 && y == 7'd44) || (x == 570 && y == 187) || (x == 7'd201 && y == 7'd555) ||
		(x == 7'd417 && y == 7'd526) || (x == 170 && y == 7'd468) || (x == 338 && y == 7'd610) ||
		(x == 7'd469 && y == 603) || (x == 577 && y == 7'd172) || (x == 7'd548 && y == 515) ||
		(x == 7'd258 && y == 7'd580) || (x == 7'd449 && y == 36) || (x == 7'd250 && y == 30) ||
		(x == 68 && y == 7'd76) || (x == 7'd330 && y == 7'd552) || (x == 608 && y == 270) ||
		(x == 7'd361 && y == 230) || (x == 7'd390 && y == 193) || (x == 7'd159 && y == 7'd374) ||
		(x == 108 && y == 7'd536) || (x == 337 && y == 7'd204) || (x == 565 && y == 7'd503) ||
		(x == 112 && y == 7'd472) || (x == 7'd452 && y == 342) || (x == 307 && y == 620) ||
		(x == 7'd504 && y == 7'd5) || (x == 7'd120 && y == 7'd83) || (x == 27 && y == 7'd434) ||
		(x == 85 && y == 7'd500) || (x == 7'd344 && y == 7'd244) || (x == 7'd19 && y == 7'd426) ||
		(x == 7'd379 && y == 613) || (x == 563 && y == 7'd256) || (x == 7'd413 && y == 7'd380) ||
		(x == 7'd19 && y == 457) || (x == 271 && y == 7'd575) || (x == 125 && y == 7'd179) ||
		(x == 178 && y == 7'd466) || (x == 7'd64 && y == 7'd348) || (x == 7'd510 && y == 7'd275) ||
		(x == 250 && y == 7'd157) || (x == 496 && y == 7'd16) || (x == 7'd510 && y == 193) ||
		(x == 7'd488 && y == 588) || (x == 417 && y == 560) || (x == 7'd622 && y == 7'd631) ||
		(x == 507 && y == 466) || (x == 153 && y == 436) || (x == 7'd497 && y == 7'd41) ||
		(x == 211 && y == 7'd18) || (x == 349 && y == 7'd632) || (x == 7'd632 && y == 181) ||
		(x == 7'd148 && y == 285) || (x == 7'd630 && y == 7'd233) || (x == 7'd197 && y == 7'd355) ||
		(x == 83 && y == 7'd299) || (x == 419 && y == 7'd437) || (x == 7'd493 && y == 7'd514) ||
		(x == 460 && y == 399) || (x == 520 && y == 223) || (x == 7'd38 && y == 269) ||
		(x == 538 && y == 7'd222) || (x == 7'd367 && y == 7'd249) || (x == 7'd409 && y == 472) ||
		(x == 7'd158 && y == 7'd380) || (x == 7'd38 && y == 7'd346) || (x == 227 && y == 7'd333) ||
		(x == 7'd463 && y == 155) || (x == 7'd367 && y == 7'd579) || (x == 310 && y == 528) ||
		(x == 7'd35 && y == 7'd531) || (x == 43 && y == 7'd491) || (x == 7'd426 && y == 7'd339) ||
		(x == 7'd191 && y == 7'd387) || (x == 308 && y == 362) || (x == 7'd69 && y == 7'd251) ||
		(x == 7'd159 && y == 7'd377) || (x == 241 && y == 300) || (x == 240 && y == 7'd470) ||
		(x == 162 && y == 7'd470) || (x == 71 && y == 7'd238) || (x == 609 && y == 343) ||
		(x == 387 && y == 407) || (x == 7'd518 && y == 7'd564) || (x == 321 && y == 7'd296) ||
		(x == 7'd49 && y == 7'd141) || (x == 316 && y == 7'd267) || (x == 298 && y == 610) ||
		(x == 112 && y == 7'd312) || (x == 7'd41 && y == 7'd527) || (x == 7'd61 && y == 7'd491) ||
		(x == 221 && y == 233) || (x == 395 && y == 164) || (x == 7'd627 && y == 7'd471) ||
		(x == 7'd285 && y == 512) || (x == 246 && y == 7'd112) || (x == 419 && y == 340) ||
		(x == 105 && y == 7'd609) || (x == 422 && y == 7'd375) || (x == 7'd204 && y == 7'd564) ||
		(x == 562 && y == 480) || (x == 7'd457 && y == 44) || (x == 7'd486 && y == 7'd260) ||
		(x == 7'd539 && y == 7'd393) || (x == 7'd200 && y == 7'd427) || (x == 488 && y == 7'd272) ||
		(x == 62 && y == 68) || (x == 7'd360 && y == 7'd299) || (x == 7'd144 && y == 161) ||
		(x == 7'd471 && y == 7'd549) || (x == 7'd283 && y == 7'd432) || (x == 7'd134 && y == 28) ||
		(x == 63 && y == 7'd172) || (x == 7'd499 && y == 7'd470) || (x == 7'd394 && y == 7'd43) ||
		(x == 7'd287 && y == 590) || (x == 37 && y == 7'd3) || (x == 281 && y == 7'd388) ||
		(x == 7'd146 && y == 7'd245) || (x == 456 && y == 7'd375) || (x == 7'd8 && y == 7'd270) ||
		(x == 7'd139 && y == 7'd627) || (x == 7'd466 && y == 7'd619) || (x == 7'd378 && y == 7'd392) ||
		(x == 5 && y == 7'd541) || (x == 7'd12 && y == 7'd112) || (x == 7'd312 && y == 7'd233) ||
		(x == 7'd533 && y == 7'd418) || (x == 7'd351 && y == 580) || (x == 7'd610 && y == 418) ||
		(x == 7'd382 && y == 7'd68) || (x == 7'd548 && y == 282) || (x == 7'd583 && y == 35) ||
		(x == 7'd483 && y == 5) || (x == 81 && y == 7'd536) || (x == 305 && y == 7'd593) ||
		(x == 7'd594 && y == 7'd433) || (x == 121 && y == 7'd469) || (x == 7'd473 && y == 7'd468) ||
		(x == 7'd387 && y == 7'd634) || (x == 7'd631 && y == 7'd458) || (x == 159 && y == 445) ||
		(x == 7'd280 && y == 7'd394) || (x == 618 && y == 7'd101) || (x == 111 && y == 7'd503) ||
		(x == 479 && y == 511) || (x == 7'd309 && y == 2) || (x == 277 && y == 637) ||
		(x == 7'd504 && y == 7'd33) || (x == 7'd255 && y == 7'd467) || (x == 7'd517 && y == 7'd556) ||
		(x == 278 && y == 7'd440) || (x == 7'd378 && y == 7'd381) || (x == 363 && y == 7'd344) ||
		(x == 130 && y == 7'd421) || (x == 7'd108 && y == 169) || (x == 485 && y == 7'd25) ||
		(x == 210 && y == 545) || (x == 621 && y == 7'd325) || (x == 576 && y == 210) ||
		(x == 22 && y == 7'd542) || (x == 618 && y == 7'd529) || (x == 7'd416 && y == 7'd27) ||
		(x == 441 && y == 7'd470) || (x == 118 && y == 7'd443) || (x == 7'd382 && y == 7'd567) ||
		(x == 7'd631 && y == 366) || (x == 7'd469 && y == 7'd373) || (x == 314 && y == 177) ||
		(x == 7'd204 && y == 7'd430) || (x == 7'd511 && y == 7'd208) || (x == 389 && y == 261) ||
		(x == 236 && y == 329) || (x == 407 && y == 131) || (x == 7'd481 && y == 262) ||
		(x == 204 && y == 7'd203) || (x == 7'd462 && y == 113) || (x == 7'd317 && y == 62) ||
		(x == 344 && y == 7'd413) || (x == 7'd500 && y == 7'd342) || (x == 497 && y == 534) ||
		(x == 7'd158 && y == 423) || (x == 7'd343 && y == 516) || (x == 447 && y == 459) ||
		(x == 7'd627 && y == 187) || (x == 555 && y == 175) || (x == 542 && y == 7'd357) ||
		(x == 616 && y == 170) || (x == 614 && y == 263) || (x == 7'd277 && y == 265) ||
		(x == 7'd639 && y == 250) || (x == 7'd130 && y == 432) || (x == 7'd84 && y == 379) ||
		(x == 221 && y == 7'd624) || (x == 407 && y == 396) || (x == 92 && y == 8) ||
		(x == 7'd527 && y == 7'd171) || (x == 7'd494 && y == 7'd476) || (x == 7'd155 && y == 235) ||
		(x == 7'd476 && y == 7'd271) || (x == 370 && y == 479) || (x == 199 && y == 179) ||
		(x == 7'd224 && y == 7'd542) || (x == 263 && y == 546) || (x == 7'd133 && y == 7'd621) ||
		(x == 500 && y == 7'd392) || (x == 526 && y == 7'd548) || (x == 7'd368 && y == 7'd435) ||
		(x == 19 && y == 7'd153) || (x == 536 && y == 7'd357) || (x == 284 && y == 7'd141) ||
		(x == 7'd391 && y == 480) || (x == 381 && y == 7'd90) || (x == 577 && y == 7'd253) ||
		(x == 7'd262 && y == 7'd544) || (x == 7'd442 && y == 7'd323) || (x == 7'd300 && y == 7'd268) ||
		(x == 340 && y == 7'd189) || (x == 7'd190 && y == 44) || (x == 568 && y == 251) ||
		(x == 233 && y == 574) || (x == 576 && y == 7'd144) || (x == 7'd402 && y == 7'd493) ||
		(x == 7'd613 && y == 7'd357) || (x == 7'd432 && y == 595) || (x == 76 && y == 7'd344) ||
		(x == 7'd197 && y == 7'd440) || (x == 7'd22 && y == 401) || (x == 7'd454 && y == 7'd399) ||
		(x == 160 && y == 7'd150) || (x == 7'd426 && y == 7'd389) || (x == 332 && y == 7'd273) ||
		(x == 7'd214 && y == 371) || (x == 7'd389 && y == 7'd437) || (x == 7'd575 && y == 7'd452) ||
		(x == 411 && y == 7'd577) || (x == 7'd164 && y == 7'd217) || (x == 7'd25 && y == 608) ||
		(x == 7'd131 && y == 7'd331) || (x == 7'd264 && y == 439) || (x == 474 && y == 560) ||
		(x == 7'd376 && y == 7'd184) || (x == 502 && y == 529) || (x == 296 && y == 7'd373) ||
		(x == 317 && y == 7'd336) || (x == 541 && y == 543) || (x == 515 && y == 7'd180) ||
		(x == 7'd373 && y == 7'd187) || (x == 7'd441 && y == 183) || (x == 235 && y == 7'd493) ||
		(x == 7'd323 && y == 7'd574) || (x == 9 && y == 7'd537) || (x == 550 && y == 570) ||
		(x == 7'd386 && y == 7'd362) || (x == 252 && y == 334) || (x == 535 && y == 524) ||
		(x == 216 && y == 510) || (x == 7'd464 && y == 7'd252) || (x == 7'd5 && y == 94) ||
		(x == 7'd137 && y == 7'd529) || (x == 200 && y == 7'd431) || (x == 7'd572 && y == 442) ||
		(x == 481 && y == 7'd511) || (x == 209 && y == 7'd414) || (x == 7'd369 && y == 7'd371) ||
		(x == 7'd581 && y == 7'd33) || (x == 7'd198 && y == 7'd166) || (x == 371 && y == 440) ||
		(x == 7'd245 && y == 274) || (x == 146 && y == 7'd619) || (x == 7'd121 && y == 7'd339) ||
		(x == 7'd290 && y == 7'd372) || (x == 7'd19 && y == 7'd51) || (x == 7'd576 && y == 7'd375) ||
		(x == 7'd463 && y == 7'd588) || (x == 7'd449 && y == 356) || (x == 314 && y == 7'd439) ||
		(x == 83 && y == 7'd259) || (x == 487 && y == 7'd151) || (x == 7'd217 && y == 270) ||
		(x == 475 && y == 416) || (x == 635 && y == 7'd56) || (x == 7'd172 && y == 187) ||
		(x == 7'd364 && y == 7'd215) || (x == 7'd252 && y == 7'd182) || (x == 7'd577 && y == 7'd303) ||
		(x == 325 && y == 7'd547) || (x == 130 && y == 7'd372) || (x == 476 && y == 7'd212) ||
		(x == 566 && y == 7'd409) || (x == 534 && y == 255) || (x == 414 && y == 149) ||
		(x == 586 && y == 7'd125) || (x == 314 && y == 526) || (x == 7'd400 && y == 7'd631) ||
		(x == 7'd394 && y == 7'd189) || (x == 364 && y == 7'd596) || (x == 279 && y == 7'd456) ||
		(x == 512 && y == 294) || (x == 307 && y == 486) || (x == 610 && y == 435) ||
		(x == 7'd364 && y == 85) || (x == 337 && y == 7'd133) || (x == 7'd579 && y == 7'd504) ||
		(x == 7'd450 && y == 7'd264) || (x == 7'd167 && y == 7'd500) || (x == 7'd625 && y == 630) ||
		(x == 7'd598 && y == 7'd481) || (x == 7'd252 && y == 7'd630) || (x == 7'd386 && y == 453) ||
		(x == 460 && y == 7'd294) || (x == 105 && y == 7'd470) || (x == 421 && y == 435) ||
		(x == 11 && y == 7'd240) || (x == 398 && y == 475) || (x == 608 && y == 172) ||
		(x == 7'd104 && y == 7'd635) || (x == 375 && y == 242) || (x == 228 && y == 190) ||
		(x == 7'd580 && y == 7'd314) || (x == 7'd582 && y == 586) || (x == 7'd241 && y == 7'd635) ||
		(x == 166 && y == 460) || (x == 7'd524 && y == 7'd595) || (x == 634 && y == 7'd547) ||
		(x == 7'd458 && y == 7'd256) || (x == 393 && y == 242) || (x == 245 && y == 593) ||
		(x == 7'd491 && y == 7'd277) || (x == 7'd522 && y == 7'd568) || (x == 623 && y == 7'd504) ||
		(x == 7'd261 && y == 613) || (x == 7'd625 && y == 7'd605) || (x == 151 && y == 622) ||
		(x == 7'd34 && y == 383) || (x == 7'd165 && y == 30) || (x == 7'd405 && y == 7'd387) ||
		(x == 7'd445 && y == 290) || (x == 175 && y == 515) || (x == 7'd266 && y == 374) ||
		(x == 7'd426 && y == 194) || (x == 7'd187 && y == 7'd385) || (x == 7'd165 && y == 230) ||
		(x == 7'd320 && y == 7'd363) || (x == 7'd304 && y == 7'd637) || (x == 577 && y == 553) ||
		(x == 414 && y == 7'd197) || (x == 7'd265 && y == 7'd335) || (x == 601 && y == 291) ||
		(x == 7'd579 && y == 7'd328) || (x == 514 && y == 570) || (x == 7'd514 && y == 7'd158) ||
		(x == 7'd619 && y == 149) || (x == 7'd188 && y == 7'd575) || (x == 7'd446 && y == 7'd325) ||
		(x == 7'd213 && y == 7'd370) || (x == 7'd293 && y == 392) || (x == 132 && y == 380) ||
		(x == 7'd76 && y == 567) || (x == 7'd602 && y == 7'd224) || (x == 424 && y == 339) ||
		(x == 8 && y == 63) || (x == 230 && y == 7'd369) || (x == 7'd353 && y == 574) ||
		(x == 563 && y == 7'd320) || (x == 165 && y == 7'd357) || (x == 7'd68 && y == 7'd253) ||
		(x == 616 && y == 244) || (x == 7'd190 && y == 155) || (x == 303 && y == 275) ||
		(x == 597 && y == 7'd622) || (x == 7'd600 && y == 7'd521) || (x == 637 && y == 7'd47) ||
		(x == 567 && y == 7'd158) || (x == 7'd220 && y == 7'd493) || (x == 7'd427 && y == 7'd318) ||
		(x == 460 && y == 7'd24) || (x == 247 && y == 361) || (x == 7'd524 && y == 390) ||
		(x == 7'd248 && y == 7'd392) || (x == 488 && y == 243) || (x == 235 && y == 7'd271) ||
		(x == 7'd451 && y == 7'd61) || (x == 7'd457 && y == 7'd414) || (x == 162 && y == 558) ||
		(x == 7'd322 && y == 7'd200) || (x == 74 && y == 7'd400) || (x == 7'd329 && y == 7'd483) ||
		(x == 155 && y == 534) || (x == 7'd189 && y == 7'd242) || (x == 228 && y == 7'd53) ||
		(x == 7'd202 && y == 7'd275) || (x == 212 && y == 7'd205) || (x == 7'd311 && y == 297) ||
		(x == 7'd585 && y == 383) || (x == 591 && y == 7'd471) || (x == 7'd495 && y == 566) ||
		(x == 190 && y == 7'd192) || (x == 7'd289 && y == 214) || (x == 7'd105 && y == 619) ||
		(x == 7'd446 && y == 7'd573) || (x == 602 && y == 227) || (x == 496 && y == 196) ||
		(x == 165 && y == 7'd581) || (x == 7'd512 && y == 483) || (x == 7'd511 && y == 7'd145) ||
		(x == 7'd639 && y == 7'd207) || (x == 7'd194 && y == 7'd284) || (x == 7'd380 && y == 7'd145) ||
		(x == 202 && y == 178) || (x == 294 && y == 7'd413) || (x == 7'd284 && y == 7'd521) ||
		(x == 7'd556 && y == 7'd137) || (x == 7'd316 && y == 156) || (x == 73 && y == 7'd256) ||
		(x == 244 && y == 7'd264) || (x == 7'd60 && y == 7'd414) || (x == 585 && y == 7'd458) ||
		(x == 520 && y == 244) || (x == 217 && y == 7'd246) || (x == 7'd325 && y == 7'd378) ||
		(x == 596 && y == 7'd214) || (x == 7'd288 && y == 7'd63) || (x == 316 && y == 285) ||
		(x == 7'd155 && y == 262) || (x == 7'd518 && y == 7'd437) || (x == 7'd486 && y == 544) ||
		(x == 183 && y == 7'd298) || (x == 241 && y == 7'd2) || (x == 196 && y == 510) ||
		(x == 7'd200 && y == 7'd285) || (x == 7'd253 && y == 620) || (x == 406 && y == 196) ||
		(x == 7'd186 && y == 7'd260) || (x == 7'd569 && y == 593) || (x == 7'd7 && y == 480) ||
		(x == 289 && y == 585) || (x == 83 && y == 7'd130) || (x == 7'd505 && y == 348) ||
		(x == 99 && y == 7'd253) || (x == 7'd185 && y == 151) || (x == 293 && y == 7'd55) ||
		(x == 501 && y == 412) || (x == 7'd636 && y == 7'd169) || (x == 7'd132 && y == 375) ||
		(x == 7'd239 && y == 316) || (x == 528 && y == 7'd395) || (x == 7'd175 && y == 370) ||
		(x == 391 && y == 433) || (x == 7'd377 && y == 7'd193) || (x == 7'd494 && y == 7'd477) ||
		(x == 7'd157 && y == 283) || (x == 7'd344 && y == 159) || (x == 7'd480 && y == 491) ||
		(x == 7'd121 && y == 7'd529) || (x == 7'd598 && y == 473) || (x == 7'd166 && y == 480) ||
		(x == 423 && y == 258) || (x == 7'd544 && y == 7'd142) || (x == 558 && y == 376) ||
		(x == 135 && y == 7'd211) || (x == 183 && y == 7'd604) || (x == 7'd172 && y == 7'd325) ||
		(x == 7'd519 && y == 63) || (x == 7'd499 && y == 571) || (x == 635 && y == 7'd178) ||
		(x == 546 && y == 7'd626) || (x == 628 && y == 7'd190) || (x == 620 && y == 480) ||
		(x == 7'd302 && y == 7'd292) || (x == 165 && y == 7'd343) || (x == 7'd400 && y == 7'd171) ||
		(x == 7'd67 && y == 7'd453) || (x == 427 && y == 7'd82) || (x == 7'd179 && y == 7'd270) ||
		(x == 584 && y == 7'd262) || (x == 7'd134 && y == 75) || (x == 7'd510 && y == 7'd205) ||
		(x == 7'd80 && y == 482) || (x == 7'd588 && y == 48) || (x == 412 && y == 324) ||
		(x == 7'd464 && y == 440) || (x == 179 && y == 7'd357) || (x == 313 && y == 405) ||
		(x == 7'd407 && y == 7'd261) || (x == 7'd261 && y == 7'd52) || (x == 483 && y == 7'd220) ||
		(x == 248 && y == 7'd612) || (x == 93 && y == 7'd271) || (x == 10 && y == 7'd93) ||
		(x == 7'd469 && y == 354) || (x == 569 && y == 7'd490) || (x == 7'd159 && y == 507) ||
		(x == 282 && y == 140) || (x == 285 && y == 7'd104) || (x == 350 && y == 7'd413) ||
		(x == 7'd250 && y == 55) || (x == 7'd481 && y == 7'd274) || (x == 7'd224 && y == 7'd143) ||
		(x == 276 && y == 589) || (x == 169 && y == 7'd55) || (x == 571 && y == 7'd532) ||
		(x == 345 && y == 256) || (x == 159 && y == 7'd56) || (x == 143 && y == 458) ||
		(x == 609 && y == 7'd345) || (x == 145 && y == 7'd531) || (x == 404 && y == 485) ||
		(x == 430 && y == 7'd311) || (x == 7'd343 && y == 7'd297) || (x == 7'd509 && y == 309) ||
		(x == 518 && y == 222) || (x == 7'd443 && y == 7'd340) || (x == 378 && y == 321) ||
		(x == 7'd174 && y == 230) || (x == 7'd102 && y == 549) || (x == 460 && y == 7'd605) ||
		(x == 7'd26 && y == 481) || (x == 7'd383 && y == 7'd225) || (x == 7'd416 && y == 7'd412) ||
		(x == 533 && y == 218) || (x == 7'd522 && y == 7'd601) || (x == 7'd382 && y == 636) ||
		(x == 7'd389 && y == 7'd283) || (x == 7'd135 && y == 222) || (x == 7'd264 && y == 7'd12) ||
		(x == 7'd607 && y == 7'd422) || (x == 139 && y == 7'd448) || (x == 588 && y == 346) ||
		(x == 225 && y == 7'd377) || (x == 7'd523 && y == 7'd497) || (x == 7'd475 && y == 7'd116) ||
		(x == 216 && y == 7'd1) || (x == 7'd452 && y == 586) || (x == 7'd421 && y == 7'd402) ||
		(x == 7'd211 && y == 311) || (x == 588 && y == 7'd271) || (x == 314 && y == 161) ||
		(x == 7'd328 && y == 7'd589) || (x == 7'd452 && y == 7'd572) || (x == 530 && y == 569) ||
		(x == 7'd185 && y == 7'd444) || (x == 7'd275 && y == 7'd271) || (x == 7'd540 && y == 579) ||
		(x == 7'd172 && y == 7'd202) || (x == 7'd145 && y == 7'd214) || (x == 7'd567 && y == 7'd147) ||
		(x == 7'd251 && y == 7'd318) || (x == 274 && y == 7'd211) || (x == 538 && y == 154) ||
		(x == 7'd573 && y == 7'd142) || (x == 529 && y == 585) || (x == 7'd318 && y == 365) ||
		(x == 7'd251 && y == 7'd157) || (x == 7'd38 && y == 513) || (x == 304 && y == 166) ||
		(x == 458 && y == 7'd297) || (x == 7'd337 && y == 7'd249) || (x == 7'd293 && y == 91) ||
		(x == 432 && y == 7'd573) || (x == 7'd160 && y == 7'd325) || (x == 7'd94 && y == 620) ||
		(x == 7'd157 && y == 7'd595) || (x == 7'd323 && y == 7'd631) || (x == 7'd307 && y == 7'd144) ||
		(x == 7'd149 && y == 52) || (x == 174 && y == 361) || (x == 35 && y == 7'd373) ||
		(x == 635 && y == 7'd308) || (x == 566 && y == 7'd85) || (x == 7'd457 && y == 371) ||
		(x == 7'd359 && y == 246) || (x == 7'd112 && y == 296) || (x == 7'd410 && y == 348) ||
		(x == 211 && y == 7'd491) || (x == 271 && y == 514) || (x == 7'd344 && y == 7'd154) ||
		(x == 619 && y == 7'd431) || (x == 7'd48 && y == 266) || (x == 7'd160 && y == 386) ||
		(x == 608 && y == 7'd532) || (x == 7'd527 && y == 19) || (x == 7'd573 && y == 527) ||
		(x == 617 && y == 7'd603) || (x == 516 && y == 185) || (x == 346 && y == 362) ||
		(x == 7'd304 && y == 282) || (x == 7'd278 && y == 7'd433) || (x == 7'd387 && y == 436) ||
		(x == 156 && y == 7'd339) || (x == 7'd238 && y == 7'd425) || (x == 145 && y == 132) ||
		(x == 7'd263 && y == 7'd460) || (x == 162 && y == 7'd625) || (x == 629 && y == 635) ||
		(x == 365 && y == 7'd154) || (x == 7'd525 && y == 7'd548) || (x == 7'd421 && y == 7'd361) ||
		(x == 7'd2 && y == 212) || (x == 7'd484 && y == 168) || (x == 7'd388 && y == 7'd137) ||
		(x == 7'd568 && y == 7'd382) || (x == 7'd213 && y == 7'd257) || (x == 115 && y == 7'd444) ||
		(x == 7'd18 && y == 372) || (x == 7'd392 && y == 277) || (x == 7'd532 && y == 510) ||
		(x == 608 && y == 7'd408) || (x == 494 && y == 7'd2) || (x == 141 && y == 173) ||
		(x == 7'd176 && y == 623) || (x == 7'd194 && y == 7'd338) || (x == 626 && y == 164) ||
		(x == 7'd144 && y == 7'd557) || (x == 7'd443 && y == 16) || (x == 7'd398 && y == 7'd188) ||
		(x == 7'd441 && y == 88) || (x == 135 && y == 209) || (x == 7'd277 && y == 601) ||
		(x == 7'd201 && y == 165) || (x == 573 && y == 7'd287) || (x == 7'd286 && y == 170) ||
		(x == 7'd625 && y == 7'd547) || (x == 7'd230 && y == 383) || (x == 362 && y == 7'd10) ||
		(x == 7'd139 && y == 325) || (x == 7'd468 && y == 455) || (x == 7'd484 && y == 7'd239) ||
		(x == 572 && y == 7'd455) || (x == 611 && y == 7'd152) || (x == 609 && y == 7'd547) ||
		(x == 7'd395 && y == 7'd237) || (x == 7'd323 && y == 7'd519) || (x == 7'd43 && y == 7'd294) ||
		(x == 7'd607 && y == 195) || (x == 7'd440 && y == 72) || (x == 550 && y == 272) ||
		(x == 7'd307 && y == 589) || (x == 258 && y == 7'd39) || (x == 7'd605 && y == 112) ||
		(x == 7'd278 && y == 226) || (x == 7'd164 && y == 7'd479) || (x == 530 && y == 341) ||
		(x == 7'd125 && y == 435) || (x == 7'd231 && y == 77) || (x == 7'd289 && y == 7'd378) ||
		(x == 415 && y == 7'd497) || (x == 7'd164 && y == 543) || (x == 7'd611 && y == 242) ||
		(x == 7'd169 && y == 7'd595) || (x == 7'd371 && y == 601) || (x == 262 && y == 7'd533) ||
		(x == 7'd296 && y == 7'd144) || (x == 7'd253 && y == 608) || (x == 7'd576 && y == 554) ||
		(x == 7'd426 && y == 7'd241) || (x == 7'd430 && y == 526) || (x == 7'd298 && y == 7'd340) ||
		(x == 179 && y == 7'd63) || (x == 111 && y == 7'd120) || (x == 7'd356 && y == 7'd285) ||
		(x == 7'd619 && y == 543) || (x == 7'd494 && y == 7'd307) || (x == 426 && y == 7'd387) ||
		(x == 7'd388 && y == 262) || (x == 7'd505 && y == 373) || (x == 7'd576 && y == 262) ||
		(x == 7'd558 && y == 4) || (x == 7'd448 && y == 186) || (x == 280 && y == 547) ||
		(x == 307 && y == 282) || (x == 7'd631 && y == 7'd600) || (x == 7'd83 && y == 7'd446) ||
		(x == 7'd124 && y == 390) || (x == 565 && y == 7'd383) || (x == 7'd27 && y == 124) ||
		(x == 444 && y == 7'd586) || (x == 7'd521 && y == 7'd216) || (x == 265 && y == 327) ||
		(x == 510 && y == 7'd328) || (x == 7'd467 && y == 7'd246) || (x == 317 && y == 219) ||
		(x == 7'd18 && y == 11) || (x == 7'd424 && y == 498) || (x == 356 && y == 7'd181) ||
		(x == 549 && y == 7'd309) || (x == 7'd62 && y == 233) || (x == 290 && y == 567) ||
		(x == 7'd391 && y == 349) || (x == 7'd362 && y == 7'd559) || (x == 7'd569 && y == 7'd212) ||
		(x == 478 && y == 208) || (x == 64 && y == 7'd322) || (x == 7'd195 && y == 7'd506) ||
		(x == 487 && y == 261) || (x == 623 && y == 7'd125) || (x == 140 && y == 7'd167) ||
		(x == 404 && y == 175) || (x == 7'd126 && y == 7'd534) || (x == 422 && y == 7'd481) ||
		(x == 7'd406 && y == 7'd140) || (x == 418 && y == 381) || (x == 7'd585 && y == 7'd403) ||
		(x == 7'd137 && y == 7'd364) || (x == 7'd241 && y == 318) || (x == 7'd581 && y == 453) ||
		(x == 207 && y == 287) || (x == 7'd133 && y == 7'd582) || (x == 183 && y == 350) ||
		(x == 489 && y == 7'd382) || (x == 615 && y == 7'd191) || (x == 7'd469 && y == 7'd617) ||
		(x == 180 && y == 7'd597) || (x == 7'd572 && y == 7'd513) || (x == 45 && y == 7'd636) ||
		(x == 412 && y == 498) || (x == 7'd602 && y == 151) || (x == 7'd467 && y == 227) ||
		(x == 7'd254 && y == 158) || (x == 7'd452 && y == 7'd251) || (x == 7'd256 && y == 471) ||
		(x == 351 && y == 7'd502) || (x == 307 && y == 7'd585) || (x == 572 && y == 506) ||
		(x == 7'd450 && y == 389) || (x == 522 && y == 7'd533) || (x == 7'd547 && y == 7'd402) ||
		(x == 7'd134 && y == 7'd477) || (x == 163 && y == 158) || (x == 7'd581 && y == 7'd523) ||
		(x == 7'd251 && y == 7'd578) || (x == 7'd551 && y == 7'd121) || (x == 275 && y == 332) ||
		(x == 7'd440 && y == 2) || (x == 7'd309 && y == 436) || (x == 327 && y == 355) ||
		(x == 7'd635 && y == 103) || (x == 557 && y == 7'd455) || (x == 443 && y == 7'd80) ||
		(x == 7'd442 && y == 310) || (x == 548 && y == 420) || (x == 202 && y == 7'd23) ||
		(x == 492 && y == 7'd269) || (x == 216 && y == 623) || (x == 7'd544 && y == 308) ||
		(x == 7'd505 && y == 7'd362) || (x == 7'd185 && y == 515) || (x == 7'd595 && y == 7'd565) ||
		(x == 636 && y == 241) || (x == 357 && y == 538) || (x == 7'd372 && y == 7'd456) ||
		(x == 7'd342 && y == 7'd7) || (x == 7'd498 && y == 7'd446) || (x == 7'd5 && y == 7'd390) ||
		(x == 7'd204 && y == 7'd489) || (x == 7'd260 && y == 343) || (x == 388 && y == 7'd612) ||
		(x == 257 && y == 7'd559) || (x == 235 && y == 7'd318) || (x == 66 && y == 7'd378) ||
		(x == 314 && y == 7'd577) || (x == 277 && y == 330) || (x == 459 && y == 617) ||
		(x == 7'd542 && y == 395) || (x == 354 && y == 410) || (x == 7'd43 && y == 7'd105) ||
		(x == 361 && y == 7'd604) || (x == 7'd306 && y == 7'd6) || (x == 225 && y == 7'd258) ||
		(x == 7'd204 && y == 385) || (x == 7'd322 && y == 7'd341) || (x == 199 && y == 7'd100) ||
		(x == 198 && y == 7'd525) || (x == 7'd202 && y == 7'd182) || (x == 178 && y == 7'd134) ||
		(x == 206 && y == 147) || (x == 7'd511 && y == 233) || (x == 7'd401 && y == 7'd319) ||
		(x == 475 && y == 597) || (x == 143 && y == 7'd264) || (x == 7'd402 && y == 7'd399) ||
		(x == 7'd514 && y == 187) || (x == 7'd467 && y == 385) || (x == 588 && y == 167) ||
		(x == 206 && y == 7'd406) || (x == 197 && y == 7'd32) || (x == 7'd283 && y == 275) ||
		(x == 7'd215 && y == 7'd504) || (x == 7'd491 && y == 7'd433) || (x == 504 && y == 7'd523) ||
		(x == 7'd379 && y == 7'd612) || (x == 7'd97 && y == 563) || (x == 7'd135 && y == 7'd518) ||
		(x == 7'd612 && y == 79) || (x == 405 && y == 480) || (x == 7'd155 && y == 7'd382) ||
		(x == 595 && y == 573) || (x == 7'd328 && y == 7'd183) || (x == 7'd360 && y == 7'd508) ||
		(x == 7'd348 && y == 387) || (x == 637 && y == 7'd455) || (x == 7'd534 && y == 7'd161) ||
		(x == 230 && y == 7'd495) || (x == 437 && y == 7'd218) || (x == 481 && y == 7'd606) ||
		(x == 497 && y == 7'd363) || (x == 7'd316 && y == 175) || (x == 333 && y == 7'd5) ||
		(x == 481 && y == 7'd323) || (x == 7'd157 && y == 266) || (x == 7'd133 && y == 7'd183) ||
		(x == 4 && y == 7'd288) || (x == 7'd272 && y == 7'd148) || (x == 7'd110 && y == 31) ||
		(x == 13 && y == 7'd38) || (x == 7'd135 && y == 363) || (x == 257 && y == 627) ||
		(x == 334 && y == 500) || (x == 7'd291 && y == 7'd1) || (x == 7'd272 && y == 583) ||
		(x == 251 && y == 7'd104) || (x == 7'd455 && y == 7'd233) || (x == 395 && y == 7'd631) ||
		(x == 268 && y == 7'd445) || (x == 134 && y == 7'd575) || (x == 163 && y == 7'd581) ||
		(x == 7'd425 && y == 7'd625) || (x == 491 && y == 183) || (x == 7'd462 && y == 180) ||
		(x == 640 && y == 499) || (x == 356 && y == 350) || (x == 389 && y == 528) ||
		(x == 7'd473 && y == 7'd18) || (x == 7'd191 && y == 7'd555) || (x == 7'd59 && y == 7'd102) ||
		(x == 7'd132 && y == 615) || (x == 254 && y == 604) || (x == 310 && y == 135) ||
		(x == 523 && y == 7'd496) || (x == 7'd13 && y == 317) || (x == 308 && y == 7'd535) ||
		(x == 67 && y == 7'd349) || (x == 7'd329 && y == 7'd253) || (x == 7'd264 && y == 7'd234) ||
		(x == 7'd282 && y == 365) || (x == 188 && y == 635) || (x == 258 && y == 7'd251) ||
		(x == 635 && y == 531) || (x == 7'd331 && y == 7'd599) || (x == 272 && y == 7'd67) ||
		(x == 7'd339 && y == 581) || (x == 125 && y == 7'd335) || (x == 7'd272 && y == 7'd18) ||
		(x == 7'd400 && y == 247) || (x == 19 && y == 7'd546) || (x == 7'd470 && y == 7'd514) ||
		(x == 195 && y == 7'd637) || (x == 546 && y == 441) || (x == 633 && y == 7'd544) ||
		(x == 7'd3 && y == 7'd516) || (x == 7'd265 && y == 7'd300) || (x == 7'd423 && y == 7'd517) ||
		(x == 7'd545 && y == 377) || (x == 589 && y == 7'd606) || (x == 7'd485 && y == 7'd555) ||
		(x == 617 && y == 7'd42) || (x == 7'd394 && y == 7'd245) || (x == 356 && y == 7'd329) ||
		(x == 555 && y == 521) || (x == 7'd200 && y == 7'd436) || (x == 7'd535 && y == 7'd157) ||
		(x == 7'd70 && y == 361) || (x == 404 && y == 209) || (x == 7'd217 && y == 441) ||
		(x == 351 && y == 7'd292) || (x == 7'd314 && y == 246) || (x == 173 && y == 234) ||
		(x == 449 && y == 135) || (x == 7'd266 && y == 7'd316) || (x == 7'd69 && y == 7'd509) ||
		(x == 7'd317 && y == 608) || (x == 7'd636 && y == 7'd251) || (x == 7'd519 && y == 7'd538) ||
		(x == 405 && y == 284) || (x == 10 && y == 7'd365) || (x == 7'd423 && y == 226) ||
		(x == 466 && y == 382) || (x == 291 && y == 7'd109) || (x == 300 && y == 426) ||
		(x == 7'd302 && y == 7'd190) || (x == 207 && y == 7'd432) || (x == 556 && y == 196) ||
		(x == 256 && y == 7'd0) || (x == 548 && y == 227) || (x == 7'd559 && y == 7'd270) ||
		(x == 7'd288 && y == 205) || (x == 268 && y == 7'd551) || (x == 270 && y == 7'd268) ||
		(x == 7'd395 && y == 7'd406) || (x == 7'd602 && y == 7'd496) || (x == 583 && y == 7'd137) ||
		(x == 7'd521 && y == 7'd239) || (x == 7'd163 && y == 294) || (x == 195 && y == 538) ||
		(x == 7'd79 && y == 7'd561) || (x == 205 && y == 195) || (x == 7'd141 && y == 7'd188) ||
		(x == 5 && y == 97) || (x == 7'd239 && y == 7'd305) || (x == 245 && y == 7'd74) ||
		(x == 453 && y == 7'd592) || (x == 7'd50 && y == 7'd482) || (x == 7'd625 && y == 7'd543) ||
		(x == 7'd243 && y == 39) || (x == 7'd299 && y == 7'd263) || (x == 7'd108 && y == 130) ||
		(x == 7'd245 && y == 592) || (x == 7'd143 && y == 7'd296) || (x == 234 && y == 7'd523) ||
		(x == 7'd290 && y == 162) || (x == 354 && y == 407) || (x == 524 && y == 7'd548) ||
		(x == 186 && y == 358) || (x == 7'd510 && y == 7'd85) || (x == 300 && y == 588) ||
		(x == 7'd477 && y == 289) || (x == 87 && y == 7'd391) || (x == 146 && y == 7'd70) ||
		(x == 224 && y == 7'd444) || (x == 7'd593 && y == 7'd601) || (x == 547 && y == 542) ||
		(x == 7'd575 && y == 7'd374) || (x == 549 && y == 7'd355) || (x == 7'd582 && y == 180) ||
		(x == 7'd438 && y == 7'd71) || (x == 7'd545 && y == 7'd15) || (x == 393 && y == 7'd390) ||
		(x == 7'd591 && y == 620) || (x == 7'd181 && y == 319) || (x == 7'd305 && y == 362) ||
		(x == 279 && y == 195) || (x == 7'd439 && y == 7'd582) || (x == 7'd7 && y == 7'd96) ||
		(x == 198 && y == 7'd188) || (x == 7'd510 && y == 7'd212) || (x == 306 && y == 364) ||
		(x == 7'd521 && y == 7'd420) || (x == 241 && y == 7'd439) || (x == 7'd167 && y == 83) ||
		(x == 7'd136 && y == 382) || (x == 7'd406 && y == 7'd284) || (x == 404 && y == 460) ||
		(x == 252 && y == 7'd88) || (x == 529 && y == 7'd289) || (x == 7'd116 && y == 608) ||
		(x == 460 && y == 433) || (x == 580 && y == 466) || (x == 575 && y == 198) ||
		(x == 7'd361 && y == 424) || (x == 7'd264 && y == 7'd223) || (x == 7'd605 && y == 7'd327) ||
		(x == 463 && y == 218) || (x == 508 && y == 7'd626) || (x == 557 && y == 7'd151) ||
		(x == 573 && y == 7'd130) || (x == 7'd162 && y == 76) || (x == 7'd619 && y == 7'd386) ||
		(x == 3 && y == 7'd235) || (x == 7'd56 && y == 605) || (x == 7'd429 && y == 473) ||
		(x == 7'd169 && y == 7'd246) || (x == 7'd278 && y == 7'd205) || (x == 479 && y == 7'd356) ||
		(x == 7'd295 && y == 264) || (x == 7'd617 && y == 7'd122) || (x == 7'd612 && y == 7'd297) ||
		(x == 71 && y == 34) || (x == 7'd37 && y == 444) || (x == 7'd383 && y == 7'd277) ||
		(x == 578 && y == 7'd348) || (x == 582 && y == 7'd542) || (x == 461 && y == 7'd184) ||
		(x == 7'd597 && y == 166) || (x == 640 && y == 408) || (x == 7'd419 && y == 386) ||
		(x == 7'd485 && y == 239) || (x == 7'd278 && y == 589) || (x == 295 && y == 7'd434) ||
		(x == 331 && y == 443) || (x == 7'd284 && y == 7'd439) || (x == 617 && y == 7'd606) ||
		(x == 7'd306 && y == 7'd424) || (x == 7'd274 && y == 7'd27) || (x == 7'd519 && y == 7'd607) ||
		(x == 7'd302 && y == 13) || (x == 160 && y == 337) || (x == 419 && y == 7'd122) ||
		(x == 7'd283 && y == 507) || (x == 625 && y == 7'd171) || (x == 7'd1 && y == 591) ||
		(x == 585 && y == 7'd134) || (x == 7'd448 && y == 604) || (x == 7'd119 && y == 6) ||
		(x == 635 && y == 7'd424) || (x == 7'd460 && y == 7'd49) || (x == 7'd443 && y == 7'd496) ||
		(x == 552 && y == 7'd196) || (x == 7'd518 && y == 7'd378) || (x == 262 && y == 7'd237) ||
		(x == 7'd355 && y == 7'd463) || (x == 7'd602 && y == 7'd500) || (x == 445 && y == 189) ||
		(x == 7'd340 && y == 7'd250) || (x == 7'd253 && y == 7'd567) || (x == 7'd154 && y == 7'd508) ||
		(x == 161 && y == 592) || (x == 7'd161 && y == 7'd402) || (x == 7'd580 && y == 7'd111) ||
		(x == 269 && y == 7'd51) || (x == 7'd427 && y == 6) || (x == 7'd378 && y == 344) ||
		(x == 391 && y == 386) || (x == 7'd552 && y == 7'd395) || (x == 7'd143 && y == 547) ||
		(x == 413 && y == 7'd111) || (x == 7'd372 && y == 7'd510) || (x == 7'd14 && y == 412) ||
		(x == 7'd397 && y == 7'd275) || (x == 257 && y == 7'd196) || (x == 7'd416 && y == 7'd273) ||
		(x == 7'd9 && y == 7'd4) || (x == 7'd442 && y == 595) || (x == 564 && y == 7'd92) ||
		(x == 7'd291 && y == 154) || (x == 108 && y == 7'd301) || (x == 7'd506 && y == 7'd273) ||
		(x == 7'd554 && y == 10) || (x == 636 && y == 7'd472) || (x == 7'd405 && y == 7'd195) ||
		(x == 7'd468 && y == 7'd217) || (x == 7'd389 && y == 7'd258) || (x == 7'd537 && y == 470) ||
		(x == 408 && y == 7'd527) || (x == 7'd321 && y == 7'd592) || (x == 7'd371 && y == 7'd254) ||
		(x == 619 && y == 7'd147) || (x == 7'd171 && y == 269) || (x == 571 && y == 7'd432) ||
		(x == 7'd318 && y == 7'd169) || (x == 229 && y == 534) || (x == 444 && y == 7'd636) ||
		(x == 7'd248 && y == 574) || (x == 7'd78 && y == 175) || (x == 7'd35 && y == 433) ||
		(x == 7'd532 && y == 7'd439) || (x == 7'd366 && y == 7'd196) || (x == 72 && y == 7'd309) ||
		(x == 193 && y == 330) || (x == 7'd337 && y == 177) || (x == 203 && y == 624) ||
		(x == 7'd585 && y == 7'd54) || (x == 213 && y == 157) || (x == 7'd434 && y == 522) ||
		(x == 7'd108 && y == 86) || (x == 7'd344 && y == 7'd348) || (x == 7'd402 && y == 7'd258) ||
		(x == 270 && y == 613) || (x == 7'd448 && y == 7'd67) || (x == 233 && y == 386) ||
		(x == 7'd396 && y == 7'd498) || (x == 7'd366 && y == 7'd39) || (x == 7'd617 && y == 7'd369) ||
		(x == 262 && y == 222) || (x == 7'd265 && y == 15) || (x == 7'd449 && y == 7'd422) ||
		(x == 7'd253 && y == 7'd554) || (x == 7'd382 && y == 7'd576) || (x == 216 && y == 7'd425) ||
		(x == 441 && y == 269) || (x == 3 && y == 7'd137) || (x == 240 && y == 577) ||
		(x == 588 && y == 7'd42) || (x == 424 && y == 7'd462) || (x == 603 && y == 129) ||
		(x == 148 && y == 139) || (x == 578 && y == 317) || (x == 240 && y == 7'd481) ||
		(x == 7'd477 && y == 7'd291) || (x == 317 && y == 7'd100) || (x == 608 && y == 7'd506) ||
		(x == 629 && y == 257) || (x == 602 && y == 7'd155) || (x == 278 && y == 7'd331) ||
		(x == 7'd96 && y == 7'd393) || (x == 161 && y == 555) || (x == 7'd424 && y == 7'd368) ||
		(x == 7'd441 && y == 140) || (x == 7'd619 && y == 7'd560) || (x == 15 && y == 7'd318) ||
		(x == 513 && y == 147) || (x == 7'd205 && y == 301) || (x == 599 && y == 7'd504) ||
		(x == 560 && y == 7'd566) || (x == 7'd614 && y == 7'd558) || (x == 7'd581 && y == 333) ||
		(x == 7'd20 && y == 361) || (x == 7'd252 && y == 7'd526) || (x == 549 && y == 239) ||
		(x == 7'd555 && y == 7'd168) || (x == 7'd551 && y == 7'd387) || (x == 7'd201 && y == 7'd479) ||
		(x == 99 && y == 7'd175) || (x == 7'd229 && y == 7'd358) || (x == 7'd31 && y == 529) ||
		(x == 7'd237 && y == 7'd426) || (x == 7'd637 && y == 562) || (x == 250 && y == 7'd221) ||
		(x == 7'd144 && y == 114) || (x == 379 && y == 7'd422) || (x == 7'd229 && y == 7'd385) ||
		(x == 503 && y == 7'd244) || (x == 7'd123 && y == 2) || (x == 7'd59 && y == 532) ||
		(x == 584 && y == 7'd376) || (x == 156 && y == 7'd326) || (x == 316 && y == 205) ||
		(x == 250 && y == 350) || (x == 67 && y == 7'd202) || (x == 7'd621 && y == 307) ||
		(x == 213 && y == 557) || (x == 398 && y == 7'd499) || (x == 7'd97 && y == 140) ||
		(x == 497 && y == 384) || (x == 118 && y == 75) || (x == 351 && y == 7'd50) ||
		(x == 453 && y == 587) || (x == 7'd497 && y == 121) || (x == 7'd209 && y == 205) ||
		(x == 366 && y == 7'd326) || (x == 7'd318 && y == 30) || (x == 7'd226 && y == 195) ||
		(x == 7'd369 && y == 7'd520) || (x == 7'd204 && y == 295) || (x == 258 && y == 7'd148) ||
		(x == 7'd487 && y == 7'd339) || (x == 7'd482 && y == 7'd237) || (x == 7'd489 && y == 460) ||
		(x == 354 && y == 316) || (x == 196 && y == 227) || (x == 7'd235 && y == 7'd583) ||
		(x == 562 && y == 7'd89) || (x == 7'd366 && y == 7'd578) || (x == 7'd508 && y == 7'd461) ||
		(x == 7'd338 && y == 7'd210) || (x == 324 && y == 7'd212) || (x == 7'd128 && y == 167) ||
		(x == 7'd98 && y == 7'd509) || (x == 7'd365 && y == 316) || (x == 461 && y == 7'd75) ||
		(x == 7'd636 && y == 45) || (x == 7'd394 && y == 114) || (x == 175 && y == 330) ||
		(x == 344 && y == 270) || (x == 7'd195 && y == 7'd441) || (x == 382 && y == 7'd261) ||
		(x == 7'd55 && y == 622) || (x == 341 && y == 518) || (x == 7'd328 && y == 320) ||
		(x == 249 && y == 129) || (x == 7'd638 && y == 7'd195) || (x == 378 && y == 241) ||
		(x == 7'd248 && y == 396) || (x == 7'd625 && y == 364) || (x == 368 && y == 7'd379) ||
		(x == 416 && y == 7'd390) || (x == 301 && y == 393) || (x == 7'd18 && y == 7'd628) ||
		(x == 7'd281 && y == 173) || (x == 7'd498 && y == 286) || (x == 7'd639 && y == 7'd461) ||
		(x == 7'd21 && y == 7'd130) || (x == 261 && y == 7'd321) || (x == 520 && y == 496) ||
		(x == 7'd219 && y == 178) || (x == 7'd491 && y == 7'd597) || (x == 7'd573 && y == 501) ||
		(x == 156 && y == 418) || (x == 7'd369 && y == 7'd601) || (x == 7'd461 && y == 145) ||
		(x == 322 && y == 7'd219) || (x == 7'd489 && y == 7'd76) || (x == 506 && y == 7'd65) ||
		(x == 7'd511 && y == 7'd212) || (x == 7'd11 && y == 203) || (x == 7'd475 && y == 205) ||
		(x == 7'd54 && y == 7'd385) || (x == 7'd158 && y == 7'd171) || (x == 401 && y == 7'd475) ||
		(x == 7'd610 && y == 547) || (x == 7'd618 && y == 7'd556) || (x == 279 && y == 133) ||
		(x == 590 && y == 7'd640) || (x == 7'd524 && y == 7'd366) || (x == 501 && y == 7'd213) ||
		(x == 7'd173 && y == 218) || (x == 176 && y == 7'd225) || (x == 471 && y == 620) ||
		(x == 561 && y == 476) || (x == 7'd532 && y == 7'd518) || (x == 623 && y == 172) ||
		(x == 117 && y == 7'd599) || (x == 604 && y == 7'd111) || (x == 158 && y == 7'd575) ||
		(x == 459 && y == 7'd347) || (x == 624 && y == 7'd57) || (x == 7'd314 && y == 335) ||
		(x == 7'd387 && y == 212) || (x == 99 && y == 7'd105) || (x == 7'd209 && y == 7'd225) ||
		(x == 7'd343 && y == 71) || (x == 585 && y == 412) || (x == 267 && y == 576) ||
		(x == 527 && y == 258) || (x == 7'd190 && y == 7'd416) || (x == 522 && y == 219) ||
		(x == 541 && y == 7'd457) || (x == 7'd436 && y == 7'd431) || (x == 7'd501 && y == 508) ||
		(x == 7'd24 && y == 7'd52) || (x == 3 && y == 7'd249) || (x == 7'd319 && y == 207) ||
		(x == 7'd538 && y == 7'd44) || (x == 7'd518 && y == 7'd282) || (x == 7'd33 && y == 618) ||
		(x == 333 && y == 216) || (x == 450 && y == 7'd302) || (x == 7'd272 && y == 7'd168) ||
		(x == 7'd204 && y == 237) || (x == 7'd414 && y == 310) || (x == 7'd443 && y == 287) ||
		(x == 276 && y == 622) || (x == 198 && y == 613) || (x == 69 && y == 7'd240) ||
		(x == 332 && y == 7'd71) || (x == 7'd65 && y == 238) || (x == 304 && y == 7'd280) ||
		(x == 198 && y == 481) || (x == 117 && y == 11) || (x == 495 && y == 397) ||
		(x == 426 && y == 595) || (x == 34 && y == 7'd148) || (x == 7'd401 && y == 7'd537) ||
		(x == 628 && y == 426) || (x == 7'd136 && y == 7'd174) || (x == 7'd395 && y == 7'd214) ||
		(x == 7'd598 && y == 7'd19) || (x == 7'd258 && y == 7'd98) || (x == 7'd348 && y == 7'd509) ||
		(x == 232 && y == 547) || (x == 7'd158 && y == 521) || (x == 7'd324 && y == 7'd294) ||
		(x == 7'd63 && y == 342) || (x == 97 && y == 7'd293) || (x == 7'd424 && y == 7'd260) ||
		(x == 588 && y == 269) || (x == 31 && y == 7'd320) || (x == 514 && y == 162) ||
		(x == 7'd589 && y == 617) || (x == 7'd569 && y == 294) || (x == 7'd94 && y == 378) ||
		(x == 7'd222 && y == 7'd549) || (x == 7'd389 && y == 7'd376) || (x == 317 && y == 7'd93) ||
		(x == 7'd12 && y == 477) || (x == 636 && y == 7'd139) || (x == 7'd506 && y == 7'd184) ||
		(x == 7'd289 && y == 7'd629) || (x == 441 && y == 7'd417) || (x == 261 && y == 316) ||
		(x == 7'd1 && y == 596) || (x == 466 && y == 7'd463) || (x == 102 && y == 7'd496) ||
		(x == 468 && y == 481) || (x == 364 && y == 593) || (x == 7'd9 && y == 622) ||
		(x == 7'd453 && y == 7'd36) || (x == 278 && y == 7'd177) || (x == 588 && y == 186) ||
		(x == 445 && y == 7'd205) || (x == 7'd94 && y == 272) || (x == 470 && y == 481) ||
		(x == 7'd149 && y == 80) || (x == 354 && y == 7'd395) || (x == 7'd386 && y == 7'd635) ||
		(x == 7'd223 && y == 7'd212) || (x == 553 && y == 7'd587) || (x == 7'd326 && y == 7'd381) ||
		(x == 370 && y == 240) || (x == 7'd240 && y == 33) || (x == 593 && y == 7'd124) ||
		(x == 7'd530 && y == 26) || (x == 7'd355 && y == 7'd550) || (x == 515 && y == 7'd437) ||
		(x == 7'd377 && y == 7'd165) || (x == 360 && y == 519) || (x == 273 && y == 7'd357) ||
		(x == 7'd332 && y == 126) || (x == 7'd467 && y == 392) || (x == 7'd356 && y == 7'd108) ||
		(x == 633 && y == 257) || (x == 7'd519 && y == 7'd155) || (x == 7'd541 && y == 613) ||
		(x == 522 && y == 251) || (x == 61 && y == 123) || (x == 7'd110 && y == 435) ||
		(x == 354 && y == 194) || (x == 7'd277 && y == 7'd465) || (x == 411 && y == 451) ||
		(x == 7'd586 && y == 132) || (x == 7'd624 && y == 94) || (x == 7'd357 && y == 548) ||
		(x == 7'd357 && y == 7'd508) || (x == 481 && y == 244) || (x == 7'd373 && y == 7'd548) ||
		(x == 7'd508 && y == 7'd532) || (x == 7'd589 && y == 105) || (x == 7'd185 && y == 7'd625) ||
		(x == 102 && y == 7'd595) || (x == 95 && y == 7'd493) || (x == 367 && y == 7'd102) ||
		(x == 247 && y == 7'd360) || (x == 592 && y == 7'd86) || (x == 7'd359 && y == 21) ||
		(x == 7'd547 && y == 264) || (x == 186 && y == 7'd66) || (x == 602 && y == 189) ||
		(x == 7'd449 && y == 133) || (x == 7'd539 && y == 636) || (x == 7'd123 && y == 405) ||
		(x == 172 && y == 7'd263) || (x == 7'd422 && y == 241) || (x == 629 && y == 7'd349) ||
		(x == 258 && y == 416) || (x == 463 && y == 7'd575) || (x == 7'd329 && y == 7'd385) ||
		(x == 550 && y == 552) || (x == 7'd329 && y == 7'd306) || (x == 634 && y == 522) ||
		(x == 7'd572 && y == 7'd627) || (x == 7'd357 && y == 7'd466) || (x == 7'd505 && y == 7'd214) ||
		(x == 356 && y == 7'd423) || (x == 376 && y == 7'd199) || (x == 130 && y == 527) ||
		(x == 391 && y == 488) || (x == 7'd295 && y == 447) || (x == 7'd86 && y == 7'd121) ||
		(x == 468 && y == 198) || (x == 7'd92 && y == 274) || (x == 7'd428 && y == 453) ||
		(x == 127 && y == 7'd459) || (x == 7'd422 && y == 136) || (x == 588 && y == 280) ||
		(x == 7'd304 && y == 439) || (x == 165 && y == 358) || (x == 624 && y == 7'd431) ||
		(x == 7'd286 && y == 515) || (x == 405 && y == 7'd617) || (x == 271 && y == 536) ||
		(x == 471 && y == 530) || (x == 7'd422 && y == 7'd627) || (x == 242 && y == 602) ||
		(x == 7'd488 && y == 381) || (x == 291 && y == 411) || (x == 7'd533 && y == 7'd155) ||
		(x == 7'd228 && y == 310) || (x == 7'd530 && y == 7'd35) || (x == 7'd154 && y == 541) ||
		(x == 7'd610 && y == 7'd303) || (x == 7'd316 && y == 297) || (x == 289 && y == 7'd45) ||
		(x == 7'd319 && y == 7'd88) || (x == 583 && y == 433) || (x == 7'd253 && y == 7'd354) ||
		(x == 7'd282 && y == 7'd436) || (x == 167 && y == 7'd561) || (x == 457 && y == 420) ||
		(x == 639 && y == 578) || (x == 287 && y == 407) || (x == 7'd407 && y == 7'd411) ||
		(x == 7'd272 && y == 7'd42) || (x == 7'd158 && y == 528) || (x == 271 && y == 460) ||
		(x == 37 && y == 7'd370) || (x == 7'd132 && y == 229) || (x == 7'd545 && y == 7'd593) ||
		(x == 7'd117 && y == 7'd124) || (x == 377 && y == 7'd276) || (x == 7'd531 && y == 7'd209) ||
		(x == 101 && y == 7'd542) || (x == 7'd575 && y == 7'd602) || (x == 395 && y == 258) ||
		(x == 7'd68 && y == 407) || (x == 7'd520 && y == 7'd169) || (x == 621 && y == 214) ||
		(x == 157 && y == 628) || (x == 114 && y == 7'd550) || (x == 564 && y == 7'd154) ||
		(x == 7'd333 && y == 7'd274) || (x == 567 && y == 7'd637) || (x == 501 && y == 177) ||
		(x == 7'd61 && y == 7'd130) || (x == 434 && y == 327) || (x == 7'd465 && y == 7'd107) ||
		(x == 7'd224 && y == 164) || (x == 415 && y == 7'd91) || (x == 7'd111 && y == 7'd412) ||
		(x == 7'd557 && y == 152) || (x == 7'd182 && y == 134) || (x == 600 && y == 458) ||
		(x == 7'd466 && y == 61) || (x == 7'd268 && y == 7'd570) || (x == 563 && y == 7'd432) ||
		(x == 285 && y == 203) || (x == 7'd623 && y == 7'd601) || (x == 7'd134 && y == 7'd537) ||
		(x == 530 && y == 437) || (x == 7'd477 && y == 7'd267) || (x == 7'd531 && y == 283) ||
		(x == 111 && y == 7'd421) || (x == 7'd77 && y == 234) || (x == 7'd600 && y == 7'd536) ||
		(x == 412 && y == 7'd94) || (x == 7'd579 && y == 7'd331) || (x == 426 && y == 7'd226) ||
		(x == 563 && y == 7'd32) || (x == 12 && y == 7'd148) || (x == 7'd346 && y == 357) ||
		(x == 499 && y == 316) || (x == 390 && y == 210) || (x == 153 && y == 7'd100) ||
		(x == 12 && y == 7'd219) || (x == 7'd391 && y == 7'd394) || (x == 7'd553 && y == 7'd363) ||
		(x == 132 && y == 572) || (x == 7'd361 && y == 7'd299) || (x == 515 && y == 640) ||
		(x == 7'd218 && y == 391) || (x == 614 && y == 554) || (x == 7'd254 && y == 26) ||
		(x == 7'd255 && y == 7'd564) || (x == 7'd41 && y == 277) || (x == 7'd273 && y == 7'd277) ||
		(x == 7'd512 && y == 250) || (x == 7'd21 && y == 389) || (x == 7'd592 && y == 444) ||
		(x == 7'd197 && y == 7'd307) || (x == 7'd392 && y == 7'd431) || (x == 7'd538 && y == 7'd608) ||
		(x == 7'd519 && y == 7'd346) || (x == 310 && y == 272) || (x == 7'd308 && y == 599) ||
		(x == 7'd582 && y == 7'd624) || (x == 615 && y == 7'd397) || (x == 279 && y == 7'd310) ||
		(x == 7'd376 && y == 318) || (x == 167 && y == 286) || (x == 7'd122 && y == 7'd333) ||
		(x == 7'd442 && y == 86) || (x == 181 && y == 218) || (x == 7'd355 && y == 462) ||
		(x == 385 && y == 7'd278) || (x == 314 && y == 286) || (x == 7'd627 && y == 7'd183) ||
		(x == 7'd312 && y == 7'd453) || (x == 7'd429 && y == 99) || (x == 7'd210 && y == 7'd557) ||
		(x == 7'd167 && y == 2) || (x == 264 && y == 7'd130) || (x == 7'd211 && y == 7'd468) ||
		(x == 7'd279 && y == 7'd253) || (x == 7'd440 && y == 504) || (x == 7'd52 && y == 7'd0) ||
		(x == 7'd415 && y == 7'd268) || (x == 7'd314 && y == 7'd129) || (x == 221 && y == 534) ||
		(x == 598 && y == 7'd177) || (x == 284 && y == 390) || (x == 7'd457 && y == 334) ||
		(x == 7'd91 && y == 7'd522) || (x == 7'd348 && y == 123) || (x == 489 && y == 524) ||
		(x == 228 && y == 7'd1) || (x == 586 && y == 312) || (x == 7'd182 && y == 7'd326) ||
		(x == 597 && y == 7'd160) || (x == 521 && y == 7'd392) || (x == 489 && y == 7'd610) ||
		(x == 7'd84 && y == 7'd514) || (x == 578 && y == 383) || (x == 182 && y == 7'd395) ||
		(x == 464 && y == 416) || (x == 133 && y == 145) || (x == 298 && y == 7'd587) ||
		(x == 7'd350 && y == 614) || (x == 7'd84 && y == 7'd87) || (x == 7'd98 && y == 619) ||
		(x == 581 && y == 7'd196) || (x == 7'd190 && y == 275) || (x == 7'd577 && y == 7'd251) ||
		(x == 7'd138 && y == 604) || (x == 432 && y == 627) || (x == 7'd555 && y == 519) ||
		(x == 198 && y == 326) || (x == 7'd191 && y == 47) || (x == 7'd178 && y == 318) ||
		(x == 7'd79 && y == 7'd494) || (x == 7'd298 && y == 129) || (x == 117 && y == 7'd456) ||
		(x == 531 && y == 7'd182) || (x == 8 && y == 7'd622) || (x == 505 && y == 586) ||
		(x == 7'd475 && y == 368) || (x == 334 && y == 256) || (x == 7'd316 && y == 90) ||
		(x == 629 && y == 189) || (x == 7'd116 && y == 552) || (x == 7'd266 && y == 7'd277) ||
		(x == 153 && y == 7'd469) || (x == 264 && y == 632) || (x == 7'd515 && y == 7'd266) ||
		(x == 574 && y == 186) || (x == 331 && y == 449) || (x == 7'd287 && y == 291) ||
		(x == 7'd147 && y == 7'd502) || (x == 7'd486 && y == 563) || (x == 443 && y == 236) ||
		(x == 7'd433 && y == 227) || (x == 7'd76 && y == 317) || (x == 334 && y == 251) ||
		(x == 493 && y == 457) || (x == 7'd93 && y == 110) || (x == 42 && y == 7'd503) ||
		(x == 7'd139 && y == 7'd441) || (x == 211 && y == 476) || (x == 7'd634 && y == 7'd192) ||
		(x == 577 && y == 7'd127) || (x == 7'd427 && y == 7'd507) || (x == 408 && y == 7'd297) ||
		(x == 413 && y == 7'd553) || (x == 7'd508 && y == 7'd569) || (x == 7'd486 && y == 161) ||
		(x == 7'd168 && y == 7'd210) || (x == 7'd448 && y == 468) || (x == 243 && y == 547) ||
		(x == 7'd628 && y == 618) || (x == 244 && y == 403) || (x == 617 && y == 460) ||
		(x == 7'd524 && y == 64) || (x == 7'd191 && y == 563) || (x == 403 && y == 165) ||
		(x == 361 && y == 568) || (x == 7'd133 && y == 7'd561) || (x == 7'd386 && y == 51) ||
		(x == 7'd392 && y == 296) || (x == 253 && y == 7'd54) || (x == 404 && y == 148) ||
		(x == 7'd597 && y == 7'd79) || (x == 7'd164 && y == 189) || (x == 7'd564 && y == 7'd432) ||
		(x == 405 && y == 7'd297) || (x == 7'd185 && y == 613) || (x == 7'd248 && y == 7'd488) ||
		(x == 7'd338 && y == 463) || (x == 7'd316 && y == 7'd529) || (x == 7'd426 && y == 7'd379) ||
		(x == 7'd551 && y == 7'd198) || (x == 7'd598 && y == 537) || (x == 335 && y == 7'd334) ||
		(x == 335 && y == 7'd464) || (x == 493 && y == 140) || (x == 7'd550 && y == 573) ||
		(x == 7'd244 && y == 7'd224) || (x == 474 && y == 7'd387) || (x == 39 && y == 7'd239) ||
		(x == 205 && y == 7'd269) || (x == 383 && y == 7'd6) || (x == 165 && y == 444) ||
		(x == 240 && y == 7'd151) || (x == 7'd613 && y == 7'd568) || (x == 7'd243 && y == 325) ||
		(x == 7'd144 && y == 492) || (x == 608 && y == 549) || (x == 7'd597 && y == 7'd505) ||
		(x == 344 && y == 7'd245) || (x == 435 && y == 263) || (x == 585 && y == 414) ||
		(x == 7'd193 && y == 7'd327) || (x == 7'd524 && y == 90) || (x == 7'd17 && y == 228) ||
		(x == 7'd58 && y == 327) || (x == 273 && y == 7'd250) || (x == 541 && y == 303) ||
		(x == 7'd223 && y == 7'd526) || (x == 625 && y == 176) || (x == 7'd404 && y == 7'd309) ||
		(x == 103 && y == 7'd341) || (x == 7'd498 && y == 7'd253) || (x == 7'd338 && y == 170) ||
		(x == 7'd621 && y == 155) || (x == 194 && y == 507) || (x == 7'd233 && y == 7'd202) ||
		(x == 7'd615 && y == 7'd403) || (x == 382 && y == 388) || (x == 7'd190 && y == 7'd90) ||
		(x == 475 && y == 307) || (x == 7'd449 && y == 7'd41) || (x == 7'd588 && y == 28) ||
		(x == 7'd435 && y == 269) || (x == 7'd509 && y == 7'd581) || (x == 7'd397 && y == 7'd370) ||
		(x == 345 && y == 151) || (x == 7'd7 && y == 7'd504) || (x == 7'd270 && y == 407) ||
		(x == 126 && y == 7'd257) || (x == 504 && y == 469) || (x == 7'd149 && y == 561) ||
		(x == 7'd365 && y == 7'd50) || (x == 7'd418 && y == 547) || (x == 424 && y == 7'd638) ||
		(x == 7'd237 && y == 7'd175) || (x == 631 && y == 7'd89) || (x == 441 && y == 202) ||
		(x == 7'd388 && y == 103) || (x == 141 && y == 7'd227) || (x == 538 && y == 548) ||
		(x == 7'd80 && y == 204) || (x == 7'd162 && y == 356) || (x == 638 && y == 618) ||
		(x == 7'd11 && y == 7'd423) || (x == 406 && y == 343) || (x == 517 && y == 481) ||
		(x == 7'd504 && y == 7'd547) || (x == 7'd394 && y == 7'd476) || (x == 7'd121 && y == 270) ||
		(x == 7'd369 && y == 7'd322) || (x == 200 && y == 7'd392) || (x == 7'd199 && y == 7'd132) ||
		(x == 215 && y == 592) || (x == 7'd508 && y == 7'd515) || (x == 326 && y == 213) ||
		(x == 429 && y == 392)) begin
			vga_r = 4'h0;
			vga_g = 4'h0;
			vga_b = 4'h0;
		end
	end
endmodule
